MACRO DFFARX1_HVT
  CLASS CORE ;
  FOREIGN DFFARX1_HVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.44 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSRHQXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9612 ;
  ANTENNAPARTIALMETALAREA 4.7986 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 21.9632 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.605 2.495 19.935 2.725 ;
      RECT 17.125 2.375 17.605 2.725 ;
      RECT 16.895 2.375 17.125 4.005 ;
      RECT 16.87 2.375 16.895 2.605 ;
      RECT 16.715 3.755 16.895 4.005 ;
      RECT 13.57 3.775 16.715 4.005 ;
      RECT 13.57 2.61 13.73 2.84 ;
      RECT 13.34 2.61 13.57 4.005 ;
      RECT 12.515 2.61 13.34 2.84 ;
      RECT 12.285 2.61 12.515 4.315 ;
      RECT 12.095 3.955 12.285 4.315 ;
      RECT 7.62 3.955 12.095 4.185 ;
      RECT 7.39 3.5 7.62 4.185 ;
      RECT 6.7 3.5 7.39 3.73 ;
      RECT 6.47 3.5 6.7 4.29 ;
      RECT 4.685 4.06 6.47 4.29 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4356 ;
  ANTENNAPARTIALMETALAREA 0.342 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4734 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.63 1.725 15.67 2.695 ;
      RECT 15.35 1.685 15.63 2.695 ;
      RECT 15.29 1.685 15.35 2.025 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.0189 ;
  ANTENNAPARTIALMETALAREA 2.3813 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.1124 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 21.565 1.37 21.57 3.195 ;
      RECT 21.34 1.37 21.565 3.205 ;
      RECT 21.275 1.37 21.34 1.6 ;
      RECT 21.335 2.965 21.34 3.205 ;
      RECT 20.2 2.975 21.335 3.205 ;
      RECT 20.905 1.26 21.275 1.6 ;
      RECT 20.015 1.37 20.905 1.6 ;
      RECT 19.86 2.975 20.2 4.17 ;
      RECT 19.405 1.26 20.015 1.6 ;
      RECT 18.13 2.975 19.86 3.205 ;
      RECT 17.845 2.975 18.13 4.01 ;
      RECT 17.79 3.19 17.845 4.01 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.4117 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4469 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.43 1.81 1.88 2.725 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.3132 ;
  ANTENNAPARTIALMETALAREA 0.3432 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2667 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.125 2.065 0.605 2.78 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.265 -0.4 22.44 0.4 ;
      RECT 17.925 -0.4 18.265 1.22 ;
      RECT 16.2 -0.4 17.925 0.4 ;
      RECT 15.86 -0.4 16.2 1.325 ;
      RECT 13.175 -0.4 15.86 0.4 ;
      RECT 12.835 -0.4 13.175 0.575 ;
      RECT 9.2 -0.4 12.835 0.4 ;
      RECT 8.86 -0.4 9.2 0.815 ;
      RECT 7.73 -0.4 8.86 0.4 ;
      RECT 7.39 -0.4 7.73 0.82 ;
      RECT 4.345 -0.4 7.39 0.4 ;
      RECT 4.005 -0.4 4.345 1.595 ;
      RECT 1.64 -0.4 4.005 0.4 ;
      RECT 1.3 -0.4 1.64 1.43 ;
      RECT 0 -0.4 1.3 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.92 4.64 22.44 5.44 ;
      RECT 20.58 3.615 20.92 5.44 ;
      RECT 19.48 4.64 20.58 5.44 ;
      RECT 19.14 3.595 19.48 5.44 ;
      RECT 16.76 4.64 19.14 5.44 ;
      RECT 16.42 4.465 16.76 5.44 ;
      RECT 15.35 4.64 16.42 5.44 ;
      RECT 15.01 4.465 15.35 5.44 ;
      RECT 13.105 4.64 15.01 5.44 ;
      RECT 12.875 3.6 13.105 5.44 ;
      RECT 7.16 4.64 12.875 5.44 ;
      RECT 6.93 3.96 7.16 5.44 ;
      RECT 4.425 4.64 6.93 5.44 ;
      RECT 4.195 3.96 4.425 5.44 ;
      RECT 1.61 4.64 4.195 5.44 ;
      RECT 1.27 3.65 1.61 5.44 ;
      RECT 0 4.64 1.27 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 22.035 1.125 22.145 1.465 ;
      RECT 21.805 0.8 22.035 1.465 ;
      RECT 20.51 0.8 21.805 1.03 ;
      RECT 20.875 1.915 21.105 2.35 ;
      RECT 16.925 1.915 20.875 2.145 ;
      RECT 20.17 0.69 20.51 1.03 ;
      RECT 19.025 0.8 20.17 1.03 ;
      RECT 18.97 0.8 19.025 1.49 ;
      RECT 18.795 0.8 18.97 1.685 ;
      RECT 18.685 1.15 18.795 1.685 ;
      RECT 17.465 1.455 18.685 1.685 ;
      RECT 17.235 0.75 17.465 1.685 ;
      RECT 17.125 0.75 17.235 1.09 ;
      RECT 16.585 1.455 16.925 2.145 ;
      RECT 16.52 1.915 16.585 2.145 ;
      RECT 16.41 1.915 16.52 2.755 ;
      RECT 16.29 1.915 16.41 3.255 ;
      RECT 16.18 2.415 16.29 3.255 ;
      RECT 16.11 3.025 16.18 3.255 ;
      RECT 15.77 3.025 16.11 3.365 ;
      RECT 15.105 3.025 15.77 3.255 ;
      RECT 15.25 1.15 15.5 1.38 ;
      RECT 15.02 0.825 15.25 1.38 ;
      RECT 14.875 2.42 15.105 3.255 ;
      RECT 13.54 0.825 15.02 1.055 ;
      RECT 14.695 2.42 14.875 2.65 ;
      RECT 14.625 1.345 14.68 1.575 ;
      RECT 14.435 1.285 14.625 1.575 ;
      RECT 14.205 1.285 14.435 3.3 ;
      RECT 12.835 1.285 14.205 1.515 ;
      RECT 14.03 3.07 14.205 3.3 ;
      RECT 13.8 3.07 14.03 3.46 ;
      RECT 13.745 1.85 13.975 2.325 ;
      RECT 11.75 2.095 13.745 2.325 ;
      RECT 12.605 1.285 12.835 1.86 ;
      RECT 12.495 1.52 12.605 1.86 ;
      RECT 11.38 3.33 12.05 3.56 ;
      RECT 11.675 2.795 11.995 3.025 ;
      RECT 11.75 0.69 11.805 0.92 ;
      RECT 11.675 0.69 11.75 2.325 ;
      RECT 11.445 0.69 11.675 3.025 ;
      RECT 10.645 0.795 11.445 1.025 ;
      RECT 10.71 2.795 11.445 3.025 ;
      RECT 11.15 3.33 11.38 3.645 ;
      RECT 10.98 1.46 11.21 2.045 ;
      RECT 8.08 3.415 11.15 3.645 ;
      RECT 9.86 1.815 10.98 2.045 ;
      RECT 10.37 2.74 10.71 3.08 ;
      RECT 10.415 0.795 10.645 1.585 ;
      RECT 10.195 1.355 10.415 1.585 ;
      RECT 9.79 0.75 10.085 0.98 ;
      RECT 9.6 2.74 9.94 3.08 ;
      RECT 9.47 1.515 9.86 2.045 ;
      RECT 9.56 0.75 9.79 1.28 ;
      RECT 8.54 2.795 9.6 3.025 ;
      RECT 7.865 1.05 9.56 1.28 ;
      RECT 8.54 1.815 9.47 2.045 ;
      RECT 8.31 1.515 8.54 3.08 ;
      RECT 8.095 1.515 8.31 1.745 ;
      RECT 7.865 3.015 8.08 3.645 ;
      RECT 7.85 1.05 7.865 3.645 ;
      RECT 7.635 1.05 7.85 3.245 ;
      RECT 6.93 1.255 7.635 1.485 ;
      RECT 6.94 3.015 7.635 3.245 ;
      RECT 7.175 1.77 7.405 2.52 ;
      RECT 5.775 1.77 7.175 2 ;
      RECT 6.82 1.2 6.93 1.54 ;
      RECT 6.59 0.655 6.82 1.54 ;
      RECT 6.235 2.235 6.755 2.465 ;
      RECT 6.42 0.655 6.59 0.885 ;
      RECT 6.005 2.235 6.235 3.675 ;
      RECT 3.47 3.445 6.005 3.675 ;
      RECT 5.665 1.445 5.775 3.215 ;
      RECT 5.545 1.39 5.665 3.215 ;
      RECT 5.325 1.39 5.545 1.73 ;
      RECT 4.415 2.985 5.545 3.215 ;
      RECT 3.015 2.115 5.31 2.345 ;
      RECT 4.185 2.595 4.415 3.215 ;
      RECT 3.86 2.595 4.185 2.825 ;
      RECT 3.24 3.03 3.47 4.41 ;
      RECT 2.54 4.17 3.24 4.41 ;
      RECT 3.005 1.225 3.015 2.345 ;
      RECT 2.98 1.225 3.005 3.91 ;
      RECT 2.775 1.17 2.98 3.91 ;
      RECT 2.64 1.17 2.775 1.51 ;
      RECT 2.5 3.045 2.54 4.41 ;
      RECT 2.27 1.93 2.5 4.41 ;
      RECT 1.07 3.045 2.27 3.275 ;
      RECT 0.87 1.2 1.07 3.275 ;
      RECT 0.84 1.145 0.87 3.275 ;
      RECT 0.53 1.145 0.84 1.485 ;
      RECT 0.73 3.045 0.84 3.275 ;
      RECT 0.445 3.045 0.73 4.195 ;
      RECT 0.39 3.375 0.445 4.195 ;
  END
END DFFARX1_HVT

MACRO SDFFX1_LVT
  CLASS CORE ;
  FOREIGN SDFFX1_LVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSRHQXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5688 ;
  ANTENNAPARTIALMETALAREA 4.0051 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 18.5235 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.91 2.61 15.14 2.95 ;
      RECT 13.93 2.665 14.91 2.895 ;
      RECT 13.7 2.25 13.93 4.235 ;
      RECT 10.47 4.005 13.7 4.235 ;
      RECT 10.43 3.01 10.47 4.235 ;
      RECT 10.42 2.71 10.43 4.235 ;
      RECT 10.345 2.66 10.42 4.235 ;
      RECT 10.24 2.405 10.345 4.235 ;
      RECT 10.115 2.405 10.24 3.24 ;
      RECT 10.09 2.63 10.115 3.24 ;
      RECT 9.51 3.01 10.09 3.24 ;
      RECT 9.28 3.01 9.51 4.405 ;
      RECT 6.82 4.175 9.28 4.405 ;
      RECT 6.59 3.445 6.82 4.405 ;
      RECT 5.895 3.445 6.59 3.675 ;
      RECT 5.665 3.445 5.895 4.41 ;
      RECT 3.99 4.18 5.665 4.41 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.3256 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.575 2.25 13.315 2.69 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.027 ;
  ANTENNAPARTIALMETALAREA 0.9159 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.4096 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.6 1.845 15.625 2.075 ;
      RECT 15.37 1.33 15.6 3.61 ;
      RECT 14.56 1.33 15.37 1.56 ;
      RECT 15.005 3.38 15.37 3.61 ;
      RECT 14.665 3.38 15.005 3.72 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.144 ;
  ANTENNAPARTIALMETALAREA 0.3877 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3303 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.85 2.06 1.4 2.765 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.216 ;
  ANTENNAPARTIALMETALAREA 0.2743 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1183 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.62 3.81 0.625 4.15 ;
      RECT 0.15 3.81 0.62 4.39 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.45 -0.4 15.84 0.4 ;
      RECT 13.11 -0.4 13.45 1.555 ;
      RECT 9.79 -0.4 13.11 0.4 ;
      RECT 9.45 -0.4 9.79 0.575 ;
      RECT 7.11 -0.4 9.45 0.4 ;
      RECT 6.77 -0.4 7.11 1.075 ;
      RECT 3.665 -0.4 6.77 0.4 ;
      RECT 3.325 -0.4 3.665 0.9 ;
      RECT 1.205 -0.4 3.325 0.4 ;
      RECT 0.865 -0.4 1.205 0.575 ;
      RECT 0 -0.4 0.865 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.66 4.64 15.84 5.44 ;
      RECT 15.32 4.465 15.66 5.44 ;
      RECT 13.655 4.64 15.32 5.44 ;
      RECT 13.315 4.465 13.655 5.44 ;
      RECT 12.345 4.64 13.315 5.44 ;
      RECT 12.005 4.465 12.345 5.44 ;
      RECT 10.01 4.64 12.005 5.44 ;
      RECT 9.78 3.64 10.01 5.44 ;
      RECT 6.355 4.64 9.78 5.44 ;
      RECT 6.125 3.915 6.355 5.44 ;
      RECT 3.66 4.64 6.125 5.44 ;
      RECT 3.32 4.465 3.66 5.44 ;
      RECT 1.195 4.64 3.32 5.44 ;
      RECT 0.855 4.465 1.195 5.44 ;
      RECT 0 4.64 0.855 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.51 0.87 15.66 1.1 ;
      RECT 15.28 0.795 15.51 1.1 ;
      RECT 14.205 0.795 15.28 1.025 ;
      RECT 14.98 1.94 15.09 2.28 ;
      RECT 14.75 1.79 14.98 2.28 ;
      RECT 12.69 1.79 14.75 2.02 ;
      RECT 14.17 0.795 14.205 1.5 ;
      RECT 13.975 0.795 14.17 1.555 ;
      RECT 13.83 1.215 13.975 1.555 ;
      RECT 13.21 2.975 13.32 3.205 ;
      RECT 12.98 2.975 13.21 3.775 ;
      RECT 12.345 2.975 12.98 3.205 ;
      RECT 11.885 3.545 12.98 3.775 ;
      RECT 12.35 1.42 12.69 2.02 ;
      RECT 12.345 1.79 12.35 2.02 ;
      RECT 12.115 1.79 12.345 3.205 ;
      RECT 12 0.72 12.19 1.06 ;
      RECT 11.85 0.72 12 1.505 ;
      RECT 11.655 2.48 11.885 3.775 ;
      RECT 11.77 0.775 11.85 1.505 ;
      RECT 10.25 1.275 11.77 1.505 ;
      RECT 11.335 1.74 11.39 1.97 ;
      RECT 10.93 1.735 11.335 1.98 ;
      RECT 11.005 0.66 11.06 1 ;
      RECT 10.72 0.66 11.005 1.035 ;
      RECT 10.7 1.735 10.93 3.58 ;
      RECT 9.91 0.805 10.72 1.035 ;
      RECT 9.53 1.75 10.7 2.015 ;
      RECT 9.68 0.805 9.91 1.27 ;
      RECT 9.045 1.04 9.68 1.27 ;
      RECT 9.295 1.75 9.53 2.12 ;
      RECT 8.815 1.04 9.045 3.225 ;
      RECT 8.645 3.605 8.985 3.945 ;
      RECT 8.29 1.04 8.815 1.27 ;
      RECT 8.22 2.995 8.815 3.225 ;
      RECT 7.28 3.715 8.645 3.945 ;
      RECT 8.35 1.5 8.58 2.71 ;
      RECT 7.87 1.5 8.35 1.73 ;
      RECT 7.74 2.48 8.35 2.71 ;
      RECT 7.28 1.96 8.11 2.19 ;
      RECT 7.64 1.07 7.87 1.73 ;
      RECT 7.51 2.48 7.74 3.48 ;
      RECT 7.53 1.07 7.64 1.41 ;
      RECT 7.05 1.31 7.28 3.945 ;
      RECT 6.31 1.31 7.05 1.54 ;
      RECT 6.05 2.975 7.05 3.205 ;
      RECT 6.465 2.255 6.78 2.485 ;
      RECT 6.235 1.775 6.465 2.485 ;
      RECT 6.15 1.2 6.31 1.54 ;
      RECT 5.005 1.775 6.235 2.005 ;
      RECT 5.97 0.63 6.15 1.54 ;
      RECT 5.92 0.63 5.97 1.485 ;
      RECT 5.615 2.24 5.955 2.58 ;
      RECT 5.81 0.63 5.92 0.97 ;
      RECT 5.43 2.35 5.615 2.58 ;
      RECT 5.2 2.35 5.43 3.845 ;
      RECT 2.84 3.615 5.2 3.845 ;
      RECT 4.97 1.3 5.005 2.005 ;
      RECT 4.74 1.3 4.97 3.27 ;
      RECT 4.665 1.3 4.74 1.64 ;
      RECT 4.32 3.04 4.74 3.27 ;
      RECT 4.28 2.005 4.51 2.38 ;
      RECT 3.98 3.04 4.32 3.38 ;
      RECT 2.625 2.005 4.28 2.235 ;
      RECT 3.4 3.04 3.98 3.27 ;
      RECT 3.39 2.525 3.4 3.27 ;
      RECT 3.17 2.47 3.39 3.27 ;
      RECT 3.05 2.47 3.17 2.81 ;
      RECT 2.61 3.615 2.84 4.345 ;
      RECT 2.395 1.195 2.625 2.735 ;
      RECT 1.885 4.115 2.61 4.345 ;
      RECT 2.1 1.195 2.395 1.425 ;
      RECT 2.345 2.505 2.395 2.735 ;
      RECT 2.115 2.505 2.345 3.825 ;
      RECT 1.885 1.77 2.15 2.11 ;
      RECT 1.81 1.77 1.885 4.345 ;
      RECT 1.655 1.825 1.81 4.345 ;
      RECT 0.52 3.22 1.655 3.45 ;
      RECT 0.465 1.21 0.52 1.55 ;
      RECT 0.465 3.165 0.52 3.505 ;
      RECT 0.235 1.21 0.465 3.505 ;
      RECT 0.18 1.21 0.235 1.55 ;
      RECT 0.18 3.165 0.235 3.505 ;
  END
END SDFFX1_LVT

MACRO DFFSRXL
  CLASS CORE ;
  FOREIGN DFFSRXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.288 ;
  ANTENNAPARTIALMETALAREA 1.7536 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.2468 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.36 4.035 11.73 4.365 ;
      RECT 8.795 4.135 11.36 4.365 ;
      RECT 8.49 4.125 8.795 4.365 ;
      RECT 6.155 4.125 8.49 4.355 ;
      RECT 6.095 4.085 6.155 4.355 ;
      RECT 5.865 4.005 6.095 4.355 ;
      RECT 5.04 4.005 5.865 4.235 ;
      RECT 4.81 4.005 5.04 4.365 ;
      RECT 4.54 4.135 4.81 4.365 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2316 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.625 1.79 6.68 2.13 ;
      RECT 6.155 1.785 6.625 2.175 ;
      RECT 6.075 1.785 6.155 2.155 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5141 ;
  ANTENNAPARTIALMETALAREA 0.7101 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1853 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.12 1.095 15.36 1.435 ;
      RECT 14.89 1.095 15.12 3.455 ;
      RECT 14.715 2.965 14.89 3.455 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 0.7408 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3708 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.555 1.095 16.685 1.435 ;
      RECT 16.345 1.095 16.555 3.23 ;
      RECT 16.33 1.205 16.345 3.23 ;
      RECT 16.325 1.205 16.33 3.58 ;
      RECT 15.99 2.965 16.325 3.58 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.3333 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.215 2.155 0.875 2.66 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2317 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0335 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.01 2.25 8.575 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.125 -0.4 17.16 0.4 ;
      RECT 15.785 -0.4 16.125 0.575 ;
      RECT 14.65 -0.4 15.785 0.4 ;
      RECT 14.31 -0.4 14.65 0.575 ;
      RECT 11.455 -0.4 14.31 0.4 ;
      RECT 11.115 -0.4 11.455 0.575 ;
      RECT 8.89 -0.4 11.115 0.4 ;
      RECT 8.55 -0.4 8.89 1.485 ;
      RECT 7.115 -0.4 8.55 0.4 ;
      RECT 6.885 -0.4 7.115 0.9 ;
      RECT 4.195 -0.4 6.885 0.4 ;
      RECT 3.855 -0.4 4.195 0.9 ;
      RECT 1.33 -0.4 3.855 0.4 ;
      RECT 0.99 -0.4 1.33 0.575 ;
      RECT 0 -0.4 0.99 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.095 4.64 17.16 5.44 ;
      RECT 15.72 4.465 16.095 5.44 ;
      RECT 13.57 4.64 15.72 5.44 ;
      RECT 13.23 3.395 13.57 5.44 ;
      RECT 12.405 4.64 13.23 5.44 ;
      RECT 12.175 3.395 12.405 5.44 ;
      RECT 11.49 3.395 12.175 3.625 ;
      RECT 5.635 4.64 12.175 5.44 ;
      RECT 11.13 3.31 11.49 3.625 ;
      RECT 10.905 3.395 11.13 3.625 ;
      RECT 10.675 3.395 10.905 3.845 ;
      RECT 8.795 3.615 10.675 3.845 ;
      RECT 8.51 3.46 8.795 3.845 ;
      RECT 8.455 3.46 8.51 3.8 ;
      RECT 5.295 4.465 5.635 5.44 ;
      RECT 4.31 4.64 5.295 5.44 ;
      RECT 3.97 4.465 4.31 5.44 ;
      RECT 1.34 4.64 3.97 5.44 ;
      RECT 0.945 4.465 1.34 5.44 ;
      RECT 0 4.64 0.945 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.6 2.22 15.92 2.56 ;
      RECT 15.58 2.22 15.6 3.915 ;
      RECT 15.37 2.275 15.58 3.915 ;
      RECT 14.475 3.685 15.37 3.915 ;
      RECT 14.415 1.17 14.66 1.51 ;
      RECT 14.415 3.505 14.475 3.915 ;
      RECT 14.32 1.17 14.415 3.915 ;
      RECT 14.245 1.225 14.32 3.915 ;
      RECT 14.185 1.225 14.245 3.735 ;
      RECT 13.95 3.395 14.185 3.735 ;
      RECT 13.725 1.825 13.955 3.165 ;
      RECT 13.605 0.98 13.855 1.32 ;
      RECT 13.145 1.825 13.725 2.055 ;
      RECT 12.01 2.935 13.725 3.165 ;
      RECT 13.515 0.63 13.605 1.32 ;
      RECT 13.375 0.63 13.515 1.265 ;
      RECT 12.275 0.63 13.375 0.86 ;
      RECT 12.915 1.09 13.145 2.055 ;
      RECT 12.715 1.09 12.915 1.32 ;
      RECT 12.135 1.89 12.475 2.23 ;
      RECT 12.255 0.63 12.275 1.235 ;
      RECT 12.045 0.63 12.255 1.29 ;
      RECT 11.065 1.89 12.135 2.12 ;
      RECT 11.915 0.95 12.045 1.29 ;
      RECT 11.78 2.615 12.01 3.165 ;
      RECT 11.295 2.615 11.78 2.845 ;
      RECT 10.955 2.56 11.295 2.9 ;
      RECT 10.835 1.25 11.065 2.12 ;
      RECT 10.415 1.25 10.835 1.48 ;
      RECT 9.545 0.72 10.705 0.95 ;
      RECT 10.185 1.25 10.415 3.36 ;
      RECT 10.115 1.25 10.185 1.535 ;
      RECT 9.775 3.13 10.185 3.36 ;
      RECT 9.885 1.195 10.115 1.535 ;
      RECT 9.545 2.43 9.87 2.77 ;
      RECT 9.315 0.72 9.545 3.125 ;
      RECT 8.035 1.745 9.315 1.975 ;
      RECT 8.075 2.895 9.315 3.125 ;
      RECT 8.02 2.895 8.075 3.8 ;
      RECT 7.805 1.37 8.035 1.975 ;
      RECT 7.845 2.895 8.02 3.835 ;
      RECT 7.575 0.74 7.935 0.97 ;
      RECT 7.735 3.46 7.845 3.835 ;
      RECT 6.555 3.605 7.735 3.835 ;
      RECT 7.345 0.74 7.575 1.365 ;
      RECT 5.67 1.135 7.345 1.365 ;
      RECT 7.26 1.635 7.3 2.795 ;
      RECT 7.245 1.635 7.26 2.8 ;
      RECT 7.07 1.635 7.245 3.375 ;
      RECT 6.92 2.46 7.07 3.375 ;
      RECT 6.87 2.565 6.92 3.375 ;
      RECT 6.785 2.905 6.87 3.375 ;
      RECT 6.1 2.905 6.785 3.135 ;
      RECT 6.325 3.545 6.555 3.835 ;
      RECT 3.72 3.545 6.325 3.775 ;
      RECT 5.87 2.54 6.1 3.135 ;
      RECT 5.64 1.12 5.67 1.46 ;
      RECT 5.41 1.12 5.64 3.135 ;
      RECT 5.33 1.12 5.41 1.46 ;
      RECT 5.09 2.905 5.41 3.135 ;
      RECT 4.935 1.84 5.165 2.205 ;
      RECT 4.045 2.905 5.09 3.26 ;
      RECT 3.585 1.975 4.935 2.205 ;
      RECT 3.815 2.51 4.045 3.26 ;
      RECT 3.49 3.545 3.72 4.365 ;
      RECT 3.355 0.955 3.585 2.965 ;
      RECT 3.14 4.135 3.49 4.365 ;
      RECT 3.03 0.955 3.355 1.24 ;
      RECT 3.055 2.735 3.355 2.965 ;
      RECT 2.895 1.77 3.125 2.225 ;
      RECT 3.055 3.48 3.11 3.82 ;
      RECT 2.825 2.735 3.055 3.82 ;
      RECT 2.69 0.9 3.03 1.24 ;
      RECT 2.43 1.995 2.895 2.225 ;
      RECT 2.77 3.48 2.825 3.82 ;
      RECT 2.43 3.045 2.505 3.405 ;
      RECT 2.23 1.49 2.43 3.405 ;
      RECT 2.275 3.98 2.33 4.32 ;
      RECT 1.99 3.81 2.275 4.32 ;
      RECT 2.215 1.435 2.23 3.405 ;
      RECT 1.845 0.745 2.225 1.05 ;
      RECT 2.2 1.435 2.215 3.3 ;
      RECT 1.89 1.435 2.2 1.775 ;
      RECT 1.555 2.96 2.2 3.3 ;
      RECT 0.52 3.81 1.99 4.04 ;
      RECT 0.465 0.815 1.845 1.045 ;
      RECT 0.465 1.43 0.52 1.77 ;
      RECT 0.29 3 0.52 4.04 ;
      RECT 0.235 0.815 0.465 1.77 ;
      RECT 0.18 3 0.29 3.34 ;
      RECT 0.18 1.43 0.235 1.77 ;
  END
END DFFSRXL

MACRO DFFSRX4
  CLASS CORE ;
  FOREIGN DFFSRX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 23.76 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9792 ;
  ANTENNAPARTIALMETALAREA 2.2933 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.7113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.18 3.995 14.52 4.335 ;
      RECT 9.025 4 14.18 4.23 ;
      RECT 8.7 4 9.025 4.335 ;
      RECT 4.86 4.105 8.7 4.335 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4614 ;
  ANTENNAPARTIALMETALAREA 0.2326 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.795 2.295 7.265 2.79 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2857 ;
  ANTENNAPARTIALMETALAREA 0.9289 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1111 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 21.565 1.82 21.64 3.22 ;
      RECT 21.335 1.475 21.565 3.22 ;
      RECT 21.26 1.42 21.335 3.22 ;
      RECT 21.255 1.42 21.26 3.195 ;
      RECT 20.86 1.42 21.255 1.82 ;
      RECT 20.9 2.855 21.255 3.195 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2857 ;
  ANTENNAPARTIALMETALAREA 0.898 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0051 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.885 1.82 22.96 3.22 ;
      RECT 22.655 1.475 22.885 3.22 ;
      RECT 22.58 1.42 22.655 3.22 ;
      RECT 22.24 1.42 22.58 1.86 ;
      RECT 22.265 2.855 22.58 3.195 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2412 ;
  ANTENNAPARTIALMETALAREA 0.2922 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.73 2.445 0.93 2.785 ;
      RECT 0.14 2.405 0.73 2.785 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.306 ;
  ANTENNAPARTIALMETALAREA 0.3329 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.7225 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.51 2.385 1.62 2.725 ;
      RECT 1.28 1.87 1.51 2.725 ;
      RECT 1.105 1.87 1.28 2.1 ;
      RECT 0.875 1.845 1.105 2.1 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 23.26 -0.4 23.76 0.4 ;
      RECT 22.92 -0.4 23.26 0.575 ;
      RECT 21.88 -0.4 22.92 0.4 ;
      RECT 21.54 -0.4 21.88 0.575 ;
      RECT 20.52 -0.4 21.54 0.4 ;
      RECT 20.18 -0.4 20.52 0.575 ;
      RECT 15.35 -0.4 20.18 0.4 ;
      RECT 15.01 -0.4 15.35 1.05 ;
      RECT 12.465 -0.4 15.01 0.4 ;
      RECT 12.125 -0.4 12.465 1.145 ;
      RECT 9.865 -0.4 12.125 0.4 ;
      RECT 9.525 -0.4 9.865 1.32 ;
      RECT 7.26 -0.4 9.525 0.4 ;
      RECT 6.92 -0.4 7.26 0.86 ;
      RECT 4.54 -0.4 6.92 0.4 ;
      RECT 4.2 -0.4 4.54 0.845 ;
      RECT 1.295 -0.4 4.2 0.4 ;
      RECT 0.955 -0.4 1.295 0.575 ;
      RECT 0 -0.4 0.955 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 23.285 4.64 23.76 5.44 ;
      RECT 22.945 4.465 23.285 5.44 ;
      RECT 21.92 4.64 22.945 5.44 ;
      RECT 21.58 4.465 21.92 5.44 ;
      RECT 20.56 4.64 21.58 5.44 ;
      RECT 20.22 4.465 20.56 5.44 ;
      RECT 17.81 4.64 20.22 5.44 ;
      RECT 17.47 3.64 17.81 5.44 ;
      RECT 15.805 4.64 17.47 5.44 ;
      RECT 15.465 2.92 15.805 5.44 ;
      RECT 13.545 4.64 15.465 5.44 ;
      RECT 13.205 4.465 13.545 5.44 ;
      RECT 12.39 4.64 13.205 5.44 ;
      RECT 12.05 4.465 12.39 5.44 ;
      RECT 9.725 4.64 12.05 5.44 ;
      RECT 9.385 4.465 9.725 5.44 ;
      RECT 4.61 4.64 9.385 5.44 ;
      RECT 4.27 4.465 4.61 5.44 ;
      RECT 1.095 4.64 4.27 5.44 ;
      RECT 0.755 4.465 1.095 5.44 ;
      RECT 0 4.64 0.755 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 23.195 2.21 23.425 3.74 ;
      RECT 20.495 3.51 23.195 3.74 ;
      RECT 20.265 1.67 20.495 3.74 ;
      RECT 19.7 1.67 20.265 1.9 ;
      RECT 19.8 3.4 20.265 3.74 ;
      RECT 19.24 2.16 19.95 2.5 ;
      RECT 19.46 3.26 19.8 4.07 ;
      RECT 19.47 0.92 19.7 1.9 ;
      RECT 19.1 1.375 19.24 3.015 ;
      RECT 19.01 1.375 19.1 3.845 ;
      RECT 18.25 1.375 19.01 1.605 ;
      RECT 18.87 2.785 19.01 3.845 ;
      RECT 18.685 0.675 18.915 1.03 ;
      RECT 18.76 3.035 18.87 3.845 ;
      RECT 18.72 1.92 18.775 2.26 ;
      RECT 16.53 3.085 18.76 3.315 ;
      RECT 18.435 1.86 18.72 2.26 ;
      RECT 17.53 0.675 18.685 0.905 ;
      RECT 16.31 1.86 18.435 2.09 ;
      RECT 17.88 1.205 18.25 1.605 ;
      RECT 16.905 1.375 17.88 1.605 ;
      RECT 17.19 0.675 17.53 1.05 ;
      RECT 16.075 0.675 17.19 0.905 ;
      RECT 16.675 1.14 16.905 1.605 ;
      RECT 16.465 1.14 16.675 1.37 ;
      RECT 16.42 3.025 16.53 3.835 ;
      RECT 16.19 2.455 16.42 3.835 ;
      RECT 16.025 1.86 16.31 2.155 ;
      RECT 15.085 2.455 16.19 2.685 ;
      RECT 15.965 0.675 16.075 1.29 ;
      RECT 13.88 1.925 16.025 2.155 ;
      RECT 15.845 0.675 15.965 1.605 ;
      RECT 15.735 0.95 15.845 1.605 ;
      RECT 14.63 1.375 15.735 1.605 ;
      RECT 15.13 4.07 15.235 4.41 ;
      RECT 14.9 3.535 15.13 4.41 ;
      RECT 15.03 2.455 15.085 3.15 ;
      RECT 14.855 2.455 15.03 3.305 ;
      RECT 8.395 3.535 14.9 3.765 ;
      RECT 14.895 4.07 14.9 4.41 ;
      RECT 14.745 2.81 14.855 3.305 ;
      RECT 12.955 3.075 14.745 3.305 ;
      RECT 14.4 0.97 14.63 1.605 ;
      RECT 14.29 0.97 14.4 1.31 ;
      RECT 13.65 0.88 13.88 2.155 ;
      RECT 13.485 0.88 13.65 1.11 ;
      RECT 13.49 1.925 13.65 2.155 ;
      RECT 13.26 1.925 13.49 2.845 ;
      RECT 13.08 1.355 13.42 1.695 ;
      RECT 11.255 1.925 13.26 2.155 ;
      RECT 11.72 1.41 13.08 1.64 ;
      RECT 12.725 2.385 12.955 3.305 ;
      RECT 12.52 2.385 12.725 2.615 ;
      RECT 11.49 0.675 11.72 1.64 ;
      RECT 10.455 0.675 11.49 0.905 ;
      RECT 11.145 1.755 11.255 3.135 ;
      RECT 11.055 1.22 11.145 3.135 ;
      RECT 11.025 1.22 11.055 3.19 ;
      RECT 10.915 1.22 11.025 1.985 ;
      RECT 10.715 2.85 11.025 3.19 ;
      RECT 10.805 1.22 10.915 1.56 ;
      RECT 10.455 2.245 10.79 2.585 ;
      RECT 10.45 0.675 10.455 2.585 ;
      RECT 10.225 0.675 10.45 2.53 ;
      RECT 8.895 2.045 10.225 2.275 ;
      RECT 8.765 1.4 9.105 1.74 ;
      RECT 8.86 2.91 9.105 3.25 ;
      RECT 7.765 0.745 8.915 0.975 ;
      RECT 8.765 2.565 8.86 3.25 ;
      RECT 8.6 1.455 8.765 1.74 ;
      RECT 8.63 2.565 8.765 3.195 ;
      RECT 8.6 2.565 8.63 2.795 ;
      RECT 8.37 1.455 8.6 2.795 ;
      RECT 8.165 3.085 8.395 3.765 ;
      RECT 8.145 2.22 8.37 2.45 ;
      RECT 7.805 3.085 8.165 3.315 ;
      RECT 7.805 1.625 7.955 1.855 ;
      RECT 7.88 3.605 7.935 3.835 ;
      RECT 7.65 3.605 7.88 3.84 ;
      RECT 7.575 1.625 7.805 3.315 ;
      RECT 7.535 0.745 7.765 1.345 ;
      RECT 3.885 3.61 7.65 3.84 ;
      RECT 6.37 3.085 7.575 3.315 ;
      RECT 5.9 1.115 7.535 1.345 ;
      RECT 6.14 2.28 6.37 3.315 ;
      RECT 5.67 1.115 5.9 3.375 ;
      RECT 5.6 1.115 5.67 1.435 ;
      RECT 4.265 3.145 5.67 3.375 ;
      RECT 5.205 1.775 5.435 2.24 ;
      RECT 3.425 1.775 5.205 2.005 ;
      RECT 4.265 2.33 4.32 2.67 ;
      RECT 4.035 2.33 4.265 3.375 ;
      RECT 3.98 2.33 4.035 2.67 ;
      RECT 3.655 3.61 3.885 4.41 ;
      RECT 2.79 4.18 3.655 4.41 ;
      RECT 3.355 0.665 3.425 2.005 ;
      RECT 3.25 0.665 3.355 2.415 ;
      RECT 3.125 0.665 3.25 3.805 ;
      RECT 3.04 0.665 3.125 0.895 ;
      RECT 3.02 2.185 3.125 3.805 ;
      RECT 2.175 1.52 2.81 1.86 ;
      RECT 2.56 3.13 2.79 4.41 ;
      RECT 2.275 0.63 2.655 1.045 ;
      RECT 2.175 3.13 2.56 3.36 ;
      RECT 2.03 3.74 2.33 4.1 ;
      RECT 0.735 0.815 2.275 1.045 ;
      RECT 1.945 1.445 2.175 3.36 ;
      RECT 0.52 3.815 2.03 4.045 ;
      RECT 1.765 1.445 1.945 1.675 ;
      RECT 1.505 3.02 1.945 3.36 ;
      RECT 0.505 0.815 0.735 1.555 ;
      RECT 0.29 3.215 0.52 4.045 ;
      RECT 0.395 1.325 0.505 1.555 ;
      RECT 0.18 3.215 0.29 3.555 ;
  END
END DFFSRX4

MACRO DFFSRX2
  CLASS CORE ;
  FOREIGN DFFSRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5328 ;
  ANTENNAPARTIALMETALAREA 1.8011 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.3846 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.17 4.035 11.665 4.365 ;
      RECT 11.005 4.085 11.17 4.365 ;
      RECT 8.525 4.135 11.005 4.365 ;
      RECT 8.295 4.125 8.525 4.365 ;
      RECT 5.9 4.125 8.295 4.355 ;
      RECT 5.67 4.005 5.9 4.355 ;
      RECT 4.845 4.005 5.67 4.235 ;
      RECT 4.615 4.005 4.845 4.365 ;
      RECT 4.345 4.135 4.615 4.365 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2268 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.085 1.77 6.625 2.19 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5865 ;
  ANTENNAPARTIALMETALAREA 0.621 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9839 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.14 1.19 15.295 1.53 ;
      RECT 14.965 1.19 15.14 3.205 ;
      RECT 14.91 1.19 14.965 3.335 ;
      RECT 14.68 2.965 14.91 3.335 ;
      RECT 14.625 3.105 14.68 3.335 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.6464 ;
  ANTENNAPARTIALMETALAREA 1.0129 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.0439 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.84 2.955 16.945 3.195 ;
      RECT 16.82 1.105 16.84 3.195 ;
      RECT 16.815 1.105 16.82 4.14 ;
      RECT 16.61 1.05 16.815 4.14 ;
      RECT 16.475 1.05 16.61 1.39 ;
      RECT 16.56 2.965 16.61 4.14 ;
      RECT 16.355 3.2 16.56 4.14 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.3782 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3038 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.565 2.115 1.18 2.73 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1944 ;
  ANTENNAPARTIALMETALAREA 0.3239 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.815 2.25 8.605 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.055 -0.4 17.16 0.4 ;
      RECT 15.715 -0.4 16.055 1.69 ;
      RECT 14.32 -0.4 15.715 0.4 ;
      RECT 13.98 -0.4 14.32 0.575 ;
      RECT 11.28 -0.4 13.98 0.4 ;
      RECT 10.94 -0.4 11.28 0.575 ;
      RECT 8.695 -0.4 10.94 0.4 ;
      RECT 8.355 -0.4 8.695 1.4 ;
      RECT 6.96 -0.4 8.355 0.4 ;
      RECT 6.73 -0.4 6.96 0.9 ;
      RECT 4 -0.4 6.73 0.4 ;
      RECT 3.66 -0.4 4 0.9 ;
      RECT 1.335 -0.4 3.66 0.4 ;
      RECT 0.995 -0.4 1.335 0.575 ;
      RECT 0 -0.4 0.995 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.875 4.64 17.16 5.44 ;
      RECT 15.535 4.09 15.875 5.44 ;
      RECT 13.295 4.64 15.535 5.44 ;
      RECT 12.955 3.56 13.295 5.44 ;
      RECT 12.21 4.64 12.955 5.44 ;
      RECT 11.98 3.485 12.21 5.44 ;
      RECT 10.71 3.485 11.98 3.715 ;
      RECT 5.44 4.64 11.98 5.44 ;
      RECT 10.48 3.485 10.71 3.845 ;
      RECT 8.64 3.615 10.48 3.845 ;
      RECT 8.3 3.505 8.64 3.845 ;
      RECT 5.1 4.465 5.44 5.44 ;
      RECT 4.115 4.64 5.1 5.44 ;
      RECT 3.775 4.465 4.115 5.44 ;
      RECT 1.28 4.64 3.775 5.44 ;
      RECT 0.94 4.465 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.75 2.145 16.255 2.375 ;
      RECT 15.52 2.145 15.75 3.83 ;
      RECT 14.38 3.6 15.52 3.83 ;
      RECT 14.34 1.225 14.38 3.95 ;
      RECT 14.15 1.17 14.34 3.95 ;
      RECT 14 1.17 14.15 1.51 ;
      RECT 14.02 3.665 14.15 3.95 ;
      RECT 13.68 3.665 14.02 4.005 ;
      RECT 13.61 1.825 13.84 3.165 ;
      RECT 12.825 1.825 13.61 2.055 ;
      RECT 12.015 2.935 13.61 3.165 ;
      RECT 13.465 0.78 13.52 1.12 ;
      RECT 13.18 0.745 13.465 1.12 ;
      RECT 12.08 0.745 13.18 0.975 ;
      RECT 12.595 1.275 12.825 2.055 ;
      RECT 12.46 1.275 12.595 1.505 ;
      RECT 11.995 1.855 12.225 2.23 ;
      RECT 11.795 0.745 12.08 1.12 ;
      RECT 11.675 2.88 12.015 3.22 ;
      RECT 10.87 1.855 11.995 2.085 ;
      RECT 11.74 0.78 11.795 1.12 ;
      RECT 11.62 2.88 11.675 3.11 ;
      RECT 11.39 2.615 11.62 3.11 ;
      RECT 10.535 2.615 11.39 2.845 ;
      RECT 10.64 1.335 10.87 2.085 ;
      RECT 10.22 1.335 10.64 1.565 ;
      RECT 9.345 0.735 10.51 0.965 ;
      RECT 9.99 1.335 10.22 3.27 ;
      RECT 9.975 1.335 9.99 1.62 ;
      RECT 9.92 3.04 9.99 3.27 ;
      RECT 9.635 1.28 9.975 1.62 ;
      RECT 9.58 3.04 9.92 3.38 ;
      RECT 9.365 2.525 9.675 2.755 ;
      RECT 9.345 1.745 9.365 2.755 ;
      RECT 9.115 0.735 9.345 3.225 ;
      RECT 7.88 1.745 9.115 1.975 ;
      RECT 7.92 2.995 9.115 3.225 ;
      RECT 7.69 2.995 7.92 3.835 ;
      RECT 7.65 1.37 7.88 1.975 ;
      RECT 7.42 0.745 7.74 0.975 ;
      RECT 7.58 3.46 7.69 3.835 ;
      RECT 6.36 3.605 7.58 3.835 ;
      RECT 7.19 0.745 7.42 1.365 ;
      RECT 7.11 2.46 7.2 2.8 ;
      RECT 5.475 1.135 7.19 1.365 ;
      RECT 6.88 1.6 7.11 3.375 ;
      RECT 6.86 2.46 6.88 3.375 ;
      RECT 6.82 2.515 6.86 3.375 ;
      RECT 6.59 2.905 6.82 3.375 ;
      RECT 5.905 2.905 6.59 3.135 ;
      RECT 6.13 3.545 6.36 3.835 ;
      RECT 3.525 3.545 6.13 3.775 ;
      RECT 5.675 2.54 5.905 3.135 ;
      RECT 5.445 1.12 5.475 1.46 ;
      RECT 5.215 1.12 5.445 3.135 ;
      RECT 5.135 1.12 5.215 1.46 ;
      RECT 4.895 2.905 5.215 3.135 ;
      RECT 4.74 1.84 4.97 2.205 ;
      RECT 3.85 2.905 4.895 3.26 ;
      RECT 3.39 1.975 4.74 2.205 ;
      RECT 3.62 2.51 3.85 3.26 ;
      RECT 3.295 3.545 3.525 4.365 ;
      RECT 3.16 0.955 3.39 2.965 ;
      RECT 2.945 4.135 3.295 4.365 ;
      RECT 2.835 0.955 3.16 1.24 ;
      RECT 2.86 2.735 3.16 2.965 ;
      RECT 2.7 1.77 2.93 2.225 ;
      RECT 2.63 2.735 2.86 3.82 ;
      RECT 2.495 0.9 2.835 1.24 ;
      RECT 2.235 1.995 2.7 2.225 ;
      RECT 2.235 3.18 2.33 3.655 ;
      RECT 2.035 1.455 2.235 3.655 ;
      RECT 1.81 3.98 2.15 4.32 ;
      RECT 1.66 0.695 2.07 1.06 ;
      RECT 2.005 1.4 2.035 3.655 ;
      RECT 1.695 1.4 2.005 1.74 ;
      RECT 1.5 3.18 2.005 3.465 ;
      RECT 0.52 3.98 1.81 4.21 ;
      RECT 0.64 0.83 1.66 1.06 ;
      RECT 0.635 0.83 0.64 1.625 ;
      RECT 0.41 0.83 0.635 1.68 ;
      RECT 0.29 3.15 0.52 4.21 ;
      RECT 0.295 1.34 0.41 1.68 ;
      RECT 0.18 3.15 0.29 3.49 ;
  END
END DFFSRX2

MACRO DFFSRX1
  CLASS CORE ;
  FOREIGN DFFSRX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3312 ;
  ANTENNAPARTIALMETALAREA 1.7474 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.2468 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.665 4.035 11.725 4.265 ;
      RECT 11.36 4.035 11.665 4.365 ;
      RECT 8.795 4.135 11.36 4.365 ;
      RECT 8.485 4.125 8.795 4.365 ;
      RECT 6.155 4.125 8.485 4.355 ;
      RECT 6.09 4.085 6.155 4.355 ;
      RECT 5.86 4.005 6.09 4.355 ;
      RECT 5.035 4.005 5.86 4.235 ;
      RECT 4.805 4.005 5.035 4.365 ;
      RECT 4.535 4.135 4.805 4.365 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2511 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0653 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.08 1.765 6.62 2.23 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.6507 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0051 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.115 1.155 15.23 1.495 ;
      RECT 15.115 3.115 15.155 3.455 ;
      RECT 14.89 1.155 15.115 3.455 ;
      RECT 14.885 1.165 14.89 3.455 ;
      RECT 14.815 2.965 14.885 3.455 ;
      RECT 14.735 2.965 14.815 3.4 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7213 ;
  ANTENNAPARTIALMETALAREA 0.7996 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5457 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.55 1.245 16.65 3.185 ;
      RECT 16.475 1.19 16.55 3.185 ;
      RECT 16.42 1.19 16.475 3.73 ;
      RECT 16.285 1.19 16.42 1.54 ;
      RECT 16.36 2.94 16.42 3.73 ;
      RECT 16.135 2.955 16.36 3.73 ;
      RECT 16.21 1.19 16.285 1.53 ;
      RECT 16.13 2.955 16.135 3.725 ;
      RECT 16.055 2.955 16.13 3.195 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2841 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2137 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.28 1.4 2.66 ;
      RECT 0.635 2.28 0.8 2.62 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.2357 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0441 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.005 2.25 8.58 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.865 -0.4 17.16 0.4 ;
      RECT 15.525 -0.4 15.865 0.575 ;
      RECT 14.51 -0.4 15.525 0.4 ;
      RECT 14.17 -0.4 14.51 0.575 ;
      RECT 11.47 -0.4 14.17 0.4 ;
      RECT 11.13 -0.4 11.47 0.575 ;
      RECT 8.885 -0.4 11.13 0.4 ;
      RECT 8.545 -0.4 8.885 1.485 ;
      RECT 7.11 -0.4 8.545 0.4 ;
      RECT 6.88 -0.4 7.11 0.9 ;
      RECT 4.19 -0.4 6.88 0.4 ;
      RECT 3.85 -0.4 4.19 0.9 ;
      RECT 1.425 -0.4 3.85 0.4 ;
      RECT 1.085 -0.4 1.425 0.575 ;
      RECT 0 -0.4 1.085 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.76 4.64 17.16 5.44 ;
      RECT 15.42 4.465 15.76 5.44 ;
      RECT 13.565 4.64 15.42 5.44 ;
      RECT 13.225 3.395 13.565 5.44 ;
      RECT 12.4 4.64 13.225 5.44 ;
      RECT 12.17 3.43 12.4 5.44 ;
      RECT 10.9 3.43 12.17 3.66 ;
      RECT 5.63 4.64 12.17 5.44 ;
      RECT 10.67 3.43 10.9 3.845 ;
      RECT 8.96 3.615 10.67 3.845 ;
      RECT 8.79 3.455 8.96 3.845 ;
      RECT 8.73 3.4 8.79 3.845 ;
      RECT 8.45 3.4 8.73 3.74 ;
      RECT 5.29 4.465 5.63 5.44 ;
      RECT 4.305 4.64 5.29 5.44 ;
      RECT 3.965 4.465 4.305 5.44 ;
      RECT 1.13 4.64 3.965 5.44 ;
      RECT 0.79 4.465 1.13 5.44 ;
      RECT 0 4.64 0.79 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.74 2.21 16.08 2.55 ;
      RECT 15.62 2.32 15.74 2.55 ;
      RECT 15.39 2.32 15.62 4.04 ;
      RECT 14.31 3.81 15.39 4.04 ;
      RECT 14.31 1.17 14.53 1.51 ;
      RECT 14.19 1.17 14.31 4.04 ;
      RECT 14.08 1.225 14.19 4.04 ;
      RECT 13.945 3.395 14.08 3.735 ;
      RECT 13.605 2.11 13.715 2.45 ;
      RECT 13.6 0.98 13.71 1.32 ;
      RECT 13.375 1.825 13.605 3.165 ;
      RECT 13.37 0.63 13.6 1.32 ;
      RECT 13.015 1.825 13.375 2.055 ;
      RECT 11.81 2.935 13.375 3.165 ;
      RECT 12.27 0.63 13.37 0.86 ;
      RECT 12.785 1.09 13.015 2.055 ;
      RECT 12.65 1.09 12.785 1.32 ;
      RECT 12.185 1.855 12.415 2.23 ;
      RECT 12.04 0.63 12.27 1.29 ;
      RECT 11.06 1.855 12.185 2.085 ;
      RECT 11.93 0.95 12.04 1.29 ;
      RECT 11.58 2.615 11.81 3.165 ;
      RECT 10.725 2.615 11.58 2.845 ;
      RECT 10.83 1.25 11.06 2.085 ;
      RECT 10.41 1.25 10.83 1.48 ;
      RECT 9.535 0.735 10.7 0.965 ;
      RECT 10.18 1.25 10.41 3.33 ;
      RECT 10.165 1.25 10.18 1.535 ;
      RECT 9.77 3.1 10.18 3.33 ;
      RECT 9.825 1.195 10.165 1.535 ;
      RECT 9.555 2.525 9.865 2.755 ;
      RECT 9.535 1.745 9.555 2.755 ;
      RECT 9.305 0.735 9.535 3.125 ;
      RECT 8.03 1.745 9.305 1.975 ;
      RECT 8.07 2.895 9.305 3.125 ;
      RECT 7.84 2.895 8.07 3.835 ;
      RECT 7.8 1.37 8.03 1.975 ;
      RECT 7.57 0.74 7.93 0.97 ;
      RECT 7.73 3.46 7.84 3.835 ;
      RECT 6.55 3.605 7.73 3.835 ;
      RECT 7.34 0.74 7.57 1.365 ;
      RECT 7.295 2.46 7.39 2.8 ;
      RECT 7.295 1.635 7.35 1.975 ;
      RECT 5.665 1.135 7.34 1.365 ;
      RECT 7.065 1.635 7.295 3.375 ;
      RECT 7.01 1.635 7.065 1.975 ;
      RECT 7.01 2.46 7.065 3.375 ;
      RECT 6.78 2.905 7.01 3.375 ;
      RECT 6.095 2.905 6.78 3.135 ;
      RECT 6.32 3.545 6.55 3.835 ;
      RECT 3.715 3.545 6.32 3.775 ;
      RECT 5.865 2.54 6.095 3.135 ;
      RECT 5.635 1.12 5.665 1.46 ;
      RECT 5.405 1.12 5.635 3.135 ;
      RECT 5.325 1.12 5.405 1.46 ;
      RECT 5.085 2.905 5.405 3.135 ;
      RECT 4.93 1.84 5.16 2.205 ;
      RECT 4.04 2.905 5.085 3.26 ;
      RECT 3.58 1.975 4.93 2.205 ;
      RECT 3.81 2.51 4.04 3.26 ;
      RECT 3.485 3.545 3.715 4.365 ;
      RECT 3.35 0.955 3.58 2.965 ;
      RECT 3.135 4.135 3.485 4.365 ;
      RECT 3.025 0.955 3.35 1.24 ;
      RECT 3.05 2.735 3.35 2.965 ;
      RECT 2.89 1.77 3.12 2.225 ;
      RECT 2.82 2.735 3.05 3.82 ;
      RECT 2.685 0.9 3.025 1.24 ;
      RECT 2.425 1.995 2.89 2.225 ;
      RECT 2.425 3.28 2.5 3.645 ;
      RECT 2.225 1.455 2.425 3.645 ;
      RECT 2.21 1.4 2.225 3.645 ;
      RECT 1.87 0.64 2.22 1.05 ;
      RECT 2.195 1.4 2.21 3.535 ;
      RECT 1.885 1.4 2.195 1.74 ;
      RECT 1.55 3.25 2.195 3.535 ;
      RECT 1.735 3.97 2.075 4.31 ;
      RECT 0.52 0.82 1.87 1.05 ;
      RECT 0.465 3.98 1.735 4.21 ;
      RECT 0.29 0.82 0.52 1.745 ;
      RECT 0.465 3.27 0.52 3.61 ;
      RECT 0.235 3.27 0.465 4.21 ;
      RECT 0.18 1.405 0.29 1.745 ;
      RECT 0.18 3.27 0.235 3.61 ;
  END
END DFFSRX1

MACRO DFFSHQXL
  CLASS CORE ;
  FOREIGN DFFSHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.2 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4968 ;
  ANTENNAPARTIALMETALAREA 2.5815 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.3049 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.005 2.19 11.305 2.53 ;
      RECT 10.965 2.19 11.005 2.635 ;
      RECT 10.855 2.22 10.965 2.635 ;
      RECT 10.625 2.22 10.855 4.175 ;
      RECT 5.415 3.945 10.625 4.175 ;
      RECT 5.185 2.66 5.415 4.175 ;
      RECT 5.065 2.66 5.185 2.945 ;
      RECT 4.835 2.405 5.065 2.945 ;
      RECT 4.165 2.555 4.835 2.945 ;
     END
  END SN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6172 ;
  ANTENNAPARTIALMETALAREA 0.9413 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.346 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.755 1.12 12.985 3.005 ;
      RECT 12.495 1.12 12.755 1.46 ;
      RECT 12.68 2.635 12.755 3.005 ;
      RECT 11.825 2.775 12.68 3.005 ;
      RECT 11.595 2.775 11.825 3.46 ;
      RECT 11.485 3.12 11.595 3.46 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.37 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.855 1.84 2.48 ;
      RECT 1.365 1.805 1.765 2.48 ;
      RECT 1.28 1.855 1.365 2.48 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2944 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.13 0.635 0.77 1.095 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.555 -0.4 13.2 0.4 ;
      RECT 11.215 -0.4 11.555 1.43 ;
      RECT 9.85 -0.4 11.215 0.4 ;
      RECT 9.51 -0.4 9.85 0.575 ;
      RECT 6.865 -0.4 9.51 0.4 ;
      RECT 6.635 -0.4 6.865 1.495 ;
      RECT 4.04 -0.4 6.635 0.4 ;
      RECT 3.7 -0.4 4.04 0.845 ;
      RECT 1.355 -0.4 3.7 0.4 ;
      RECT 1.015 -0.4 1.355 0.575 ;
      RECT 0 -0.4 1.015 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.545 4.64 13.2 5.44 ;
      RECT 12.205 3.32 12.545 5.44 ;
      RECT 11.215 4.64 12.205 5.44 ;
      RECT 10.875 4.465 11.215 5.44 ;
      RECT 9.835 4.64 10.875 5.44 ;
      RECT 9.495 4.465 9.835 5.44 ;
      RECT 6.66 4.64 9.495 5.44 ;
      RECT 6.295 4.465 6.66 5.44 ;
      RECT 4.95 4.64 6.295 5.44 ;
      RECT 4.01 4.14 4.95 5.44 ;
      RECT 1.45 4.64 4.01 5.44 ;
      RECT 1.11 4.465 1.45 5.44 ;
      RECT 0 4.64 1.11 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.44 2.165 12.445 2.45 ;
      RECT 12.215 1.725 12.44 2.45 ;
      RECT 12.21 1.725 12.215 2.395 ;
      RECT 10.605 1.725 12.21 1.955 ;
      RECT 10.49 0.805 10.605 1.955 ;
      RECT 10.375 0.695 10.49 1.955 ;
      RECT 10.135 0.695 10.375 1.04 ;
      RECT 10.14 2.64 10.345 3.15 ;
      RECT 10.115 1.29 10.14 3.15 ;
      RECT 9.56 0.81 10.135 1.04 ;
      RECT 9.91 1.29 10.115 2.87 ;
      RECT 9.25 2.64 9.91 2.87 ;
      RECT 9.33 0.81 9.56 2.265 ;
      RECT 8.485 0.81 9.33 1.04 ;
      RECT 8.79 2.035 9.33 2.265 ;
      RECT 9.02 2.64 9.25 3 ;
      RECT 8.33 1.485 8.9 1.715 ;
      RECT 6.725 3.44 8.865 3.67 ;
      RECT 8.56 2.035 8.79 3.19 ;
      RECT 7.92 2.96 8.56 3.19 ;
      RECT 8.145 0.755 8.485 1.095 ;
      RECT 8.1 1.485 8.33 2.445 ;
      RECT 7.71 2.215 8.1 2.445 ;
      RECT 7.615 1.105 7.725 1.445 ;
      RECT 7.48 2.215 7.71 2.58 ;
      RECT 7.385 1.105 7.615 1.965 ;
      RECT 7.235 2.96 7.41 3.19 ;
      RECT 7.235 1.735 7.385 1.965 ;
      RECT 7.005 1.735 7.235 3.19 ;
      RECT 6.495 1.87 6.725 3.67 ;
      RECT 6.395 1.87 6.495 2.1 ;
      RECT 6.375 3.395 6.495 3.67 ;
      RECT 6.165 1.35 6.395 2.1 ;
      RECT 5.645 3.395 6.375 3.625 ;
      RECT 5.935 2.33 6.26 2.67 ;
      RECT 6.065 1.35 6.165 1.58 ;
      RECT 5.835 0.675 6.065 1.58 ;
      RECT 5.92 1.81 5.935 2.67 ;
      RECT 5.705 1.81 5.92 2.615 ;
      RECT 5.5 0.675 5.835 0.905 ;
      RECT 5.55 1.81 5.705 2.04 ;
      RECT 5.32 1.335 5.55 2.04 ;
      RECT 4.96 1.335 5.32 1.995 ;
      RECT 4.625 0.775 5.065 1.005 ;
      RECT 3.935 1.765 4.96 1.995 ;
      RECT 4.32 3.34 4.66 3.68 ;
      RECT 4.395 0.775 4.625 1.365 ;
      RECT 2.99 1.135 4.395 1.365 ;
      RECT 3.935 3.34 4.32 3.57 ;
      RECT 3.705 1.765 3.935 3.57 ;
      RECT 3.315 1.885 3.705 2.115 ;
      RECT 3.245 2.36 3.475 3.635 ;
      RECT 2.985 2.36 3.245 2.59 ;
      RECT 2.775 3.405 3.245 3.635 ;
      RECT 2.34 2.87 3.015 3.1 ;
      RECT 2.985 1.015 2.99 1.365 ;
      RECT 2.755 1.015 2.985 2.59 ;
      RECT 2.435 3.405 2.775 3.745 ;
      RECT 2.675 1.015 2.755 1.3 ;
      RECT 2.335 0.96 2.675 1.3 ;
      RECT 2.11 1.715 2.34 3.1 ;
      RECT 0.89 2.87 2.11 3.1 ;
      RECT 0.59 2.87 0.89 3.49 ;
      RECT 0.59 1.345 0.645 1.685 ;
      RECT 0.55 1.345 0.59 3.49 ;
      RECT 0.36 1.345 0.55 3.1 ;
      RECT 0.305 1.345 0.36 1.685 ;
  END
END DFFSHQXL

MACRO DFFSHQX4
  CLASS CORE ;
  FOREIGN DFFSHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 18.48 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSHQXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.6884 ;
  ANTENNAPARTIALMETALAREA 3.6466 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 16.854 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.715 2.25 16.94 2.48 ;
      RECT 16.38 2.25 16.715 2.565 ;
      RECT 15.055 2.335 16.38 2.565 ;
      RECT 15.01 2.255 15.055 2.565 ;
      RECT 14.78 2.255 15.01 4.235 ;
      RECT 14.64 2.255 14.78 2.485 ;
      RECT 14.66 3.755 14.78 4.235 ;
      RECT 10.045 4.005 14.66 4.235 ;
      RECT 9.815 3.53 10.045 4.235 ;
      RECT 5.645 3.53 9.815 3.76 ;
      RECT 5.645 2.965 5.725 3.195 ;
      RECT 5.415 2.9 5.645 3.76 ;
      RECT 4.43 2.9 5.415 3.13 ;
     END
  END SN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.1228 ;
  ANTENNAPARTIALMETALAREA 2.7092 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.4569 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.28 0.8 18.3 1.29 ;
      RECT 18.05 0.8 18.28 3.185 ;
      RECT 17.96 0.8 18.05 1.495 ;
      RECT 17.68 2.955 18.05 3.185 ;
      RECT 15.74 1.265 17.96 1.495 ;
      RECT 17.3 2.94 17.68 4.34 ;
      RECT 17.08 2.985 17.3 4.03 ;
      RECT 17.02 2.985 17.08 3.22 ;
      RECT 15.98 2.985 17.02 3.215 ;
      RECT 15.9 2.985 15.98 3.22 ;
      RECT 15.56 2.985 15.9 3.925 ;
      RECT 15.505 1.055 15.74 1.495 ;
      RECT 15.4 1.055 15.505 1.395 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2988 ;
  ANTENNAPARTIALMETALAREA 0.2475 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.375 1.955 2.875 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.4428 ;
  ANTENNAPARTIALMETALAREA 0.2755 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 1.82 1.18 2.545 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 17.02 -0.4 18.48 0.4 ;
      RECT 16.68 -0.4 17.02 0.955 ;
      RECT 14.25 -0.4 16.68 0.4 ;
      RECT 12.97 -0.4 14.25 0.575 ;
      RECT 8.82 -0.4 12.97 0.4 ;
      RECT 8.48 -0.4 8.82 1.28 ;
      RECT 7.375 -0.4 8.48 0.4 ;
      RECT 7.035 -0.4 7.375 1.395 ;
      RECT 4.085 -0.4 7.035 0.4 ;
      RECT 3.745 -0.4 4.085 0.575 ;
      RECT 1.52 -0.4 3.745 0.4 ;
      RECT 1.18 -0.4 1.52 0.575 ;
      RECT 0 -0.4 1.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.215 4.64 18.48 5.44 ;
      RECT 17.985 3.48 18.215 5.44 ;
      RECT 16.66 4.64 17.985 5.44 ;
      RECT 16.32 3.48 16.66 5.44 ;
      RECT 15.1 4.64 16.32 5.44 ;
      RECT 14.76 4.465 15.1 5.44 ;
      RECT 13.63 4.64 14.76 5.44 ;
      RECT 13.29 4.465 13.63 5.44 ;
      RECT 8.95 4.64 13.29 5.44 ;
      RECT 8.61 4.465 8.95 5.44 ;
      RECT 7.425 4.64 8.61 5.44 ;
      RECT 7.085 4.465 7.425 5.44 ;
      RECT 5.96 4.64 7.085 5.44 ;
      RECT 5.62 4.465 5.96 5.44 ;
      RECT 4.44 4.64 5.62 5.44 ;
      RECT 4.1 4.465 4.44 5.44 ;
      RECT 1.73 4.64 4.1 5.44 ;
      RECT 1.39 4.465 1.73 5.44 ;
      RECT 0 4.64 1.39 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 17.71 2.205 17.82 2.545 ;
      RECT 17.48 1.78 17.71 2.545 ;
      RECT 16.08 1.78 17.48 2.01 ;
      RECT 15.68 1.78 16.08 2.065 ;
      RECT 15.015 1.78 15.68 2.01 ;
      RECT 14.785 0.865 15.015 2.01 ;
      RECT 12.205 0.865 14.785 1.095 ;
      RECT 14.31 3 14.42 3.34 ;
      RECT 14.08 1.545 14.31 3.34 ;
      RECT 13.26 1.545 14.08 1.775 ;
      RECT 13.705 2.25 13.815 2.59 ;
      RECT 13.475 2.25 13.705 3.775 ;
      RECT 12.205 3.545 13.475 3.775 ;
      RECT 12.92 1.37 13.26 1.775 ;
      RECT 12.885 1.54 12.92 1.775 ;
      RECT 12.6 1.54 12.885 2.345 ;
      RECT 12.545 2.005 12.6 2.345 ;
      RECT 11.975 0.865 12.205 3.775 ;
      RECT 11.7 0.865 11.975 1.095 ;
      RECT 10.42 3.545 11.975 3.775 ;
      RECT 11.59 0.865 11.7 1.41 ;
      RECT 11.36 0.725 11.59 1.41 ;
      RECT 10.88 3.07 11.52 3.3 ;
      RECT 10.26 0.725 11.36 0.955 ;
      RECT 10.88 1.2 10.98 1.54 ;
      RECT 10.65 1.2 10.88 3.3 ;
      RECT 10.64 1.2 10.65 1.745 ;
      RECT 7.845 3.07 10.65 3.3 ;
      RECT 9.54 1.515 10.64 1.745 ;
      RECT 10.03 0.725 10.26 1.28 ;
      RECT 9.92 0.94 10.03 1.28 ;
      RECT 7.585 1.975 10.025 2.205 ;
      RECT 9.2 1.1 9.54 1.745 ;
      RECT 9.255 3.995 9.485 4.405 ;
      RECT 3.495 3.995 9.255 4.225 ;
      RECT 8.1 1.515 9.2 1.745 ;
      RECT 7.815 1.11 8.1 1.745 ;
      RECT 7.76 1.11 7.815 1.45 ;
      RECT 7.355 1.725 7.585 3.155 ;
      RECT 6.585 1.725 7.355 1.955 ;
      RECT 6.465 2.925 7.355 3.155 ;
      RECT 5.635 2.26 7.12 2.49 ;
      RECT 6.355 0.775 6.585 1.955 ;
      RECT 4.85 0.775 6.355 1.005 ;
      RECT 5.565 1.3 5.635 2.665 ;
      RECT 5.405 1.245 5.565 2.665 ;
      RECT 5.225 1.245 5.405 1.585 ;
      RECT 3.865 2.435 5.405 2.665 ;
      RECT 3.2 1.975 5.175 2.205 ;
      RECT 4.915 3.365 5.145 3.76 ;
      RECT 3.865 3.365 4.915 3.595 ;
      RECT 4.62 0.775 4.85 1.705 ;
      RECT 3.485 1.475 4.62 1.705 ;
      RECT 3.635 2.435 3.865 3.595 ;
      RECT 3.21 3.995 3.495 4.235 ;
      RECT 3.255 0.635 3.485 1.705 ;
      RECT 3.075 0.635 3.255 0.865 ;
      RECT 2.735 4.005 3.21 4.235 ;
      RECT 3.02 1.975 3.2 3.715 ;
      RECT 2.97 1.175 3.02 3.715 ;
      RECT 2.79 1.175 2.97 2.205 ;
      RECT 2.5 1.175 2.79 1.405 ;
      RECT 2.505 3.605 2.735 4.235 ;
      RECT 2.415 3.605 2.505 3.835 ;
      RECT 2.185 1.74 2.415 3.835 ;
      RECT 0.955 3.605 2.185 3.835 ;
      RECT 0.615 3 0.955 3.94 ;
      RECT 0.57 1.18 0.76 1.52 ;
      RECT 0.57 3 0.615 3.23 ;
      RECT 0.42 1.18 0.57 3.23 ;
      RECT 0.34 1.235 0.42 3.23 ;
  END
END DFFSHQX4

MACRO DFFSHQX2
  CLASS CORE ;
  FOREIGN DFFSHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSHQXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9396 ;
  ANTENNAPARTIALMETALAREA 4.2354 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 19.0747 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.16 2.11 15.215 2.45 ;
      RECT 14.93 2.11 15.16 3.755 ;
      RECT 14.875 2.11 14.93 2.45 ;
      RECT 12.755 3.525 14.93 3.755 ;
      RECT 12.55 2.175 12.78 2.515 ;
      RECT 12.55 3.5 12.755 3.755 ;
      RECT 12.44 2.175 12.55 3.755 ;
      RECT 12.41 2.23 12.44 3.755 ;
      RECT 12.32 2.23 12.41 4.305 ;
      RECT 12.18 3.525 12.32 4.305 ;
      RECT 8.36 4.075 12.18 4.305 ;
      RECT 8.13 3.655 8.36 4.305 ;
      RECT 8.06 3.655 8.13 4.085 ;
      RECT 7.12 3.655 8.06 3.885 ;
      RECT 6.93 3.655 7.12 4.085 ;
      RECT 6.7 3.655 6.93 4.365 ;
      RECT 5.145 4.135 6.7 4.365 ;
      RECT 5.065 2.455 5.145 4.365 ;
      RECT 4.915 2.405 5.065 4.365 ;
      RECT 4.115 2.405 4.915 2.685 ;
      RECT 3.83 2.405 4.115 2.78 ;
      RECT 3.775 2.44 3.83 2.78 ;
     END
  END SN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4 ;
  ANTENNAPARTIALMETALAREA 0.8729 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9909 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.415 1.315 14.645 3.08 ;
      RECT 14.21 1.315 14.415 1.545 ;
      RECT 14.075 2.85 14.415 3.08 ;
      RECT 13.87 1.205 14.21 1.545 ;
      RECT 13.74 2.85 14.075 3.19 ;
      RECT 13.415 2.85 13.74 3.195 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.4341 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.6271 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.055 1.82 1.475 2.755 ;
      RECT 0.875 1.845 1.055 2.075 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.2293 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.475 3.805 0.675 4.235 ;
      RECT 0.215 3.805 0.475 4.315 ;
      RECT 0.19 3.805 0.215 4.235 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.49 -0.4 15.84 0.4 ;
      RECT 15.15 -0.4 15.49 1.51 ;
      RECT 12.41 -0.4 15.15 0.4 ;
      RECT 12.07 -0.4 12.41 0.575 ;
      RECT 8.285 -0.4 12.07 0.4 ;
      RECT 7.945 -0.4 8.285 1.39 ;
      RECT 6.79 -0.4 7.945 0.4 ;
      RECT 6.56 -0.4 6.79 1.37 ;
      RECT 3.865 -0.4 6.56 0.4 ;
      RECT 3.525 -0.4 3.865 0.96 ;
      RECT 1.28 -0.4 3.525 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.515 4.64 15.84 5.44 ;
      RECT 14.175 4.085 14.515 5.44 ;
      RECT 13.015 4.64 14.175 5.44 ;
      RECT 12.675 4.035 13.015 5.44 ;
      RECT 7.75 4.64 12.675 5.44 ;
      RECT 7.41 4.17 7.75 5.44 ;
      RECT 4.545 4.64 7.41 5.44 ;
      RECT 3.735 4.14 4.545 5.44 ;
      RECT 1.31 4.64 3.735 5.44 ;
      RECT 0.97 4.465 1.31 5.44 ;
      RECT 0 4.64 0.97 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.725 2.04 14.065 2.38 ;
      RECT 13.25 2.04 13.725 2.27 ;
      RECT 13.02 0.865 13.25 2.27 ;
      RECT 10.475 0.865 13.02 1.095 ;
      RECT 11.72 2.125 11.95 3.745 ;
      RECT 11.645 2.125 11.72 2.355 ;
      RECT 11.43 3.515 11.72 3.745 ;
      RECT 11.645 1.46 11.7 1.8 ;
      RECT 11.415 1.46 11.645 2.355 ;
      RECT 10.475 2.815 11.485 3.045 ;
      RECT 11.36 1.46 11.415 1.8 ;
      RECT 11.4 2.06 11.415 2.355 ;
      RECT 11.06 2.06 11.4 2.4 ;
      RECT 10.315 0.865 10.475 3.845 ;
      RECT 10.245 0.795 10.315 3.845 ;
      RECT 10.085 0.795 10.245 1.6 ;
      RECT 8.89 3.615 10.245 3.845 ;
      RECT 8.985 0.795 10.085 1.025 ;
      RECT 9.755 3.135 10.01 3.365 ;
      RECT 9.705 1.625 9.755 3.365 ;
      RECT 9.525 1.28 9.705 3.365 ;
      RECT 9.365 1.28 9.525 1.86 ;
      RECT 6.695 3.135 9.525 3.365 ;
      RECT 7.565 1.63 9.365 1.86 ;
      RECT 6.465 2.09 9.285 2.32 ;
      RECT 8.755 0.795 8.985 1.28 ;
      RECT 8.645 0.94 8.755 1.28 ;
      RECT 7.335 1.115 7.565 1.86 ;
      RECT 7.225 1.115 7.335 1.455 ;
      RECT 6.235 1.75 6.465 3.845 ;
      RECT 6.09 1.75 6.235 1.98 ;
      RECT 5.845 3.56 6.235 3.845 ;
      RECT 5.99 1.41 6.09 1.98 ;
      RECT 5.86 0.675 5.99 1.98 ;
      RECT 5.75 2.24 5.98 2.875 ;
      RECT 5.76 0.675 5.86 1.64 ;
      RECT 5.505 3.56 5.845 3.9 ;
      RECT 5.345 0.675 5.76 0.905 ;
      RECT 5.62 2.24 5.75 2.47 ;
      RECT 5.39 1.875 5.62 2.47 ;
      RECT 5.245 1.875 5.39 2.105 ;
      RECT 5.015 1.415 5.245 2.105 ;
      RECT 4.905 1.415 5.015 1.885 ;
      RECT 4.665 0.72 5.005 1.06 ;
      RECT 3.44 1.655 4.905 1.885 ;
      RECT 4.545 0.83 4.665 1.06 ;
      RECT 4.315 0.83 4.545 1.42 ;
      RECT 4.18 3.3 4.52 3.64 ;
      RECT 2.62 1.19 4.315 1.42 ;
      RECT 3.385 3.355 4.18 3.585 ;
      RECT 3.385 1.655 3.44 2.51 ;
      RECT 3.21 1.655 3.385 3.585 ;
      RECT 3.155 2.17 3.21 3.585 ;
      RECT 3.1 2.17 3.155 2.51 ;
      RECT 2.12 3.96 2.975 4.19 ;
      RECT 2.39 1.19 2.62 3.57 ;
      RECT 2.35 1.19 2.39 1.585 ;
      RECT 2.35 3.135 2.39 3.57 ;
      RECT 2.14 1.355 2.35 1.585 ;
      RECT 2.12 1.835 2.155 2.205 ;
      RECT 1.89 1.835 2.12 4.19 ;
      RECT 0.615 3.245 1.89 3.475 ;
      RECT 0.375 3.135 0.615 3.475 ;
      RECT 0.375 1.455 0.56 1.795 ;
      RECT 0.145 1.455 0.375 3.475 ;
  END
END DFFSHQX2

MACRO DFFSHQX1
  CLASS CORE ;
  FOREIGN DFFSHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.2 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSHQXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5652 ;
  ANTENNAPARTIALMETALAREA 2.7007 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 12.0522 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.435 1.845 11.665 2.1 ;
      RECT 11.305 1.87 11.435 2.1 ;
      RECT 11.075 1.87 11.305 2.45 ;
      RECT 10.965 2.11 11.075 2.45 ;
      RECT 10.855 2.22 10.965 2.45 ;
      RECT 10.625 2.22 10.855 4.175 ;
      RECT 5.415 3.945 10.625 4.175 ;
      RECT 5.185 2.66 5.415 4.175 ;
      RECT 5.065 2.66 5.185 2.945 ;
      RECT 4.835 2.405 5.065 2.945 ;
      RECT 4.165 2.555 4.835 2.945 ;
     END
  END SN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.934 ;
  ANTENNAPARTIALMETALAREA 0.9889 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5474 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.755 0.855 12.985 3.005 ;
      RECT 12.68 0.855 12.755 1.285 ;
      RECT 12.68 2.635 12.755 3.005 ;
      RECT 12.55 0.855 12.68 1.22 ;
      RECT 11.825 2.775 12.68 3.005 ;
      RECT 11.595 2.775 11.825 3.44 ;
      RECT 11.485 3.1 11.595 3.44 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3472 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.22 1.82 1.84 2.38 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.198 ;
  ANTENNAPARTIALMETALAREA 0.2812 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1872 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.675 1.18 3.22 ;
      RECT 0.605 2.675 0.8 3.055 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.595 -0.4 13.2 0.4 ;
      RECT 11.175 -0.4 11.595 1.01 ;
      RECT 9.85 -0.4 11.175 0.4 ;
      RECT 9.51 -0.4 9.85 0.575 ;
      RECT 6.865 -0.4 9.51 0.4 ;
      RECT 6.635 -0.4 6.865 1.28 ;
      RECT 4.04 -0.4 6.635 0.4 ;
      RECT 3.7 -0.4 4.04 0.845 ;
      RECT 1.28 -0.4 3.7 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.545 4.64 13.2 5.44 ;
      RECT 12.205 3.32 12.545 5.44 ;
      RECT 11.24 4.64 12.205 5.44 ;
      RECT 10.9 4.465 11.24 5.44 ;
      RECT 9.835 4.64 10.9 5.44 ;
      RECT 9.495 4.465 9.835 5.44 ;
      RECT 6.66 4.64 9.495 5.44 ;
      RECT 6.295 4.465 6.66 5.44 ;
      RECT 4.95 4.64 6.295 5.44 ;
      RECT 4.01 4.14 4.95 5.44 ;
      RECT 1.1 4.64 4.01 5.44 ;
      RECT 0.76 4.465 1.1 5.44 ;
      RECT 0 4.64 0.76 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.26 2.165 12.42 2.395 ;
      RECT 12.03 1.285 12.26 2.395 ;
      RECT 10.605 1.285 12.03 1.515 ;
      RECT 10.49 0.805 10.605 1.515 ;
      RECT 10.375 0.695 10.49 1.515 ;
      RECT 10.155 2.64 10.385 3.15 ;
      RECT 10.135 0.695 10.375 1.035 ;
      RECT 10.14 2.64 10.155 2.87 ;
      RECT 9.91 1.32 10.14 2.87 ;
      RECT 9.38 0.805 10.135 1.035 ;
      RECT 9.25 2.64 9.91 2.87 ;
      RECT 9.15 0.805 9.38 2.265 ;
      RECT 9.02 2.64 9.25 3 ;
      RECT 8.665 0.805 9.15 1.035 ;
      RECT 8.79 2.035 9.15 2.265 ;
      RECT 8.33 1.45 8.9 1.68 ;
      RECT 6.725 3.44 8.865 3.67 ;
      RECT 8.56 2.035 8.79 3.19 ;
      RECT 8.43 0.805 8.665 1.22 ;
      RECT 7.92 2.96 8.56 3.19 ;
      RECT 8.025 0.99 8.43 1.22 ;
      RECT 8.1 1.45 8.33 2.445 ;
      RECT 7.71 2.215 8.1 2.445 ;
      RECT 7.48 2.215 7.71 2.58 ;
      RECT 7.53 1.08 7.64 1.42 ;
      RECT 7.3 1.08 7.53 1.835 ;
      RECT 7.235 2.96 7.455 3.19 ;
      RECT 7.235 1.605 7.3 1.835 ;
      RECT 7.005 1.605 7.235 3.19 ;
      RECT 6.495 1.595 6.725 3.67 ;
      RECT 6.395 1.595 6.495 1.825 ;
      RECT 6.375 3.385 6.495 3.67 ;
      RECT 6.165 1.35 6.395 1.825 ;
      RECT 5.685 3.385 6.375 3.615 ;
      RECT 5.935 2.355 6.26 2.585 ;
      RECT 6.065 1.35 6.165 1.58 ;
      RECT 5.835 0.675 6.065 1.58 ;
      RECT 5.705 1.81 5.935 2.585 ;
      RECT 5.5 0.675 5.835 0.905 ;
      RECT 5.55 1.81 5.705 2.04 ;
      RECT 5.32 1.335 5.55 2.04 ;
      RECT 4.96 1.335 5.32 1.995 ;
      RECT 4.625 0.775 5.065 1.005 ;
      RECT 3.935 1.765 4.96 1.995 ;
      RECT 3.935 3.395 4.66 3.625 ;
      RECT 4.395 0.775 4.625 1.365 ;
      RECT 2.99 1.135 4.395 1.365 ;
      RECT 3.705 1.765 3.935 3.625 ;
      RECT 3.315 1.845 3.705 2.075 ;
      RECT 3.245 2.365 3.475 3.89 ;
      RECT 2.985 2.365 3.245 2.595 ;
      RECT 2.385 3.66 3.245 3.89 ;
      RECT 2.985 0.855 2.99 1.365 ;
      RECT 2.755 0.855 2.985 2.595 ;
      RECT 2.345 2.995 2.965 3.225 ;
      RECT 2.335 0.855 2.755 1.085 ;
      RECT 2.115 1.775 2.345 3.425 ;
      RECT 1.82 3.195 2.115 3.425 ;
      RECT 1.59 3.195 1.82 3.87 ;
      RECT 0.52 3.64 1.59 3.87 ;
      RECT 0.37 3.32 0.52 3.87 ;
      RECT 0.37 1.385 0.465 1.755 ;
      RECT 0.14 1.385 0.37 3.87 ;
  END
END DFFSHQX1

MACRO DFFSXL
  CLASS CORE ;
  FOREIGN DFFSXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.54 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.2091 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9752 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.38 3.9 9.79 4.41 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 1.217 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.6657 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.46 0.87 11.69 3.97 ;
      RECT 10.945 0.87 11.46 1.1 ;
      RECT 11.1 3.74 11.46 3.97 ;
      RECT 11.005 3.74 11.1 4.21 ;
      RECT 10.76 3.74 11.005 4.315 ;
      RECT 10.605 0.755 10.945 1.1 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 0.5847 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.325 3.09 12.36 3.43 ;
      RECT 12.095 1.25 12.325 3.43 ;
      RECT 11.96 1.25 12.095 1.59 ;
      RECT 12.02 3.09 12.095 3.43 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.205 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.425 1.205 1.835 1.705 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2879 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.03 2.965 1.105 3.195 ;
      RECT 0.8 2.48 1.03 3.195 ;
      RECT 0.605 2.48 0.8 2.82 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.165 -0.4 12.54 0.4 ;
      RECT 11.825 -0.4 12.165 0.575 ;
      RECT 10.22 -0.4 11.825 0.4 ;
      RECT 9.88 -0.4 10.22 1.095 ;
      RECT 8.56 -0.4 9.88 0.4 ;
      RECT 8.22 -0.4 8.56 0.575 ;
      RECT 6.165 -0.4 8.22 0.4 ;
      RECT 5.935 -0.4 6.165 1.01 ;
      RECT 4.04 -0.4 5.935 0.4 ;
      RECT 3.7 -0.4 4.04 1.09 ;
      RECT 1.535 -0.4 3.7 0.4 ;
      RECT 1.195 -0.4 1.535 0.575 ;
      RECT 0 -0.4 1.195 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.36 4.64 12.54 5.44 ;
      RECT 12.305 4.465 12.36 5.44 ;
      RECT 12.075 4.41 12.305 5.44 ;
      RECT 12.02 4.465 12.075 5.44 ;
      RECT 10.38 4.64 12.02 5.44 ;
      RECT 10.04 3.17 10.38 5.44 ;
      RECT 8.93 4.64 10.04 5.44 ;
      RECT 8.59 4.08 8.93 5.44 ;
      RECT 6.42 4.64 8.59 5.44 ;
      RECT 6.08 4.135 6.42 5.44 ;
      RECT 5.16 4.64 6.08 5.44 ;
      RECT 4.82 4.135 5.16 5.44 ;
      RECT 3.76 4.64 4.82 5.44 ;
      RECT 3.42 4.465 3.76 5.44 ;
      RECT 1.3 4.64 3.42 5.44 ;
      RECT 0.96 4.465 1.3 5.44 ;
      RECT 0 4.64 0.96 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 11.1 2.11 11.225 2.45 ;
      RECT 10.985 1.57 11.1 3.51 ;
      RECT 10.87 1.46 10.985 3.51 ;
      RECT 10.645 1.46 10.87 1.8 ;
      RECT 10.76 3.17 10.87 3.51 ;
      RECT 9.66 1.985 10.37 2.325 ;
      RECT 9.43 1.455 9.66 3.51 ;
      RECT 7.88 1.455 9.43 1.685 ;
      RECT 9.32 3.17 9.43 3.51 ;
      RECT 8.39 2.41 9.2 2.75 ;
      RECT 8.16 1.915 8.39 3.21 ;
      RECT 7.325 1.915 8.16 2.145 ;
      RECT 7.74 2.98 8.16 3.21 ;
      RECT 6.84 2.5 7.93 2.73 ;
      RECT 7.4 2.98 7.74 3.32 ;
      RECT 7.26 3.93 7.37 4.27 ;
      RECT 7.095 1.47 7.325 2.145 ;
      RECT 7.03 3.675 7.26 4.27 ;
      RECT 5.73 3.675 7.03 3.905 ;
      RECT 6.61 1.24 6.84 3.33 ;
      RECT 5.705 1.24 6.61 1.47 ;
      RECT 5.92 3.1 6.61 3.33 ;
      RECT 5.245 2.165 6.375 2.505 ;
      RECT 5.58 3.1 5.92 3.44 ;
      RECT 5.39 3.675 5.73 3.945 ;
      RECT 5.475 0.78 5.705 1.47 ;
      RECT 5.385 0.78 5.475 1.01 ;
      RECT 2.88 3.675 5.39 3.905 ;
      RECT 5.04 0.63 5.385 1.01 ;
      RECT 5.015 1.46 5.245 3.235 ;
      RECT 4.27 0.63 5.04 0.86 ;
      RECT 4.56 3.005 5.015 3.235 ;
      RECT 4.62 2.43 4.73 2.77 ;
      RECT 4.39 2.18 4.62 2.77 ;
      RECT 4.22 3.005 4.56 3.44 ;
      RECT 2.91 2.18 4.39 2.41 ;
      RECT 3.6 3.005 4.22 3.235 ;
      RECT 3.37 2.64 3.6 3.235 ;
      RECT 3.26 2.64 3.37 2.98 ;
      RECT 2.9 0.76 2.91 2.41 ;
      RECT 2.67 0.75 2.9 3.24 ;
      RECT 2.54 3.675 2.88 4.14 ;
      RECT 2.515 0.75 2.67 1.09 ;
      RECT 2.6 3.01 2.67 3.24 ;
      RECT 2.26 3.01 2.6 3.35 ;
      RECT 1.905 3.675 2.54 3.905 ;
      RECT 2.095 1.85 2.435 2.19 ;
      RECT 1.905 1.96 2.095 2.19 ;
      RECT 1.655 1.96 1.905 3.905 ;
      RECT 0.53 1.96 1.655 2.19 ;
      RECT 0.54 3.45 1.655 3.68 ;
      RECT 0.2 3.22 0.54 3.68 ;
      RECT 0.3 1.19 0.53 2.19 ;
      RECT 0.19 1.19 0.3 1.53 ;
  END
END DFFSXL

MACRO DFFSX4
  CLASS CORE ;
  FOREIGN DFFSX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 18.48 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9288 ;
  ANTENNAPARTIALMETALAREA 0.3168 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3144 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.26 4.05 5.14 4.41 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.62 ;
  ANTENNAPARTIALMETALAREA 1.033 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5881 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.21 1.82 16.36 3.22 ;
      RECT 16.06 1.26 16.21 3.22 ;
      RECT 15.98 0.855 16.06 3.22 ;
      RECT 15.72 0.855 15.98 1.665 ;
      RECT 15.6 2.78 15.98 3.12 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5984 ;
  ANTENNAPARTIALMETALAREA 1.3754 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4802 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.96 1.82 18.34 3.22 ;
      RECT 17.5 1.82 17.96 2.05 ;
      RECT 17.325 2.985 17.96 3.215 ;
      RECT 17.27 0.855 17.5 2.05 ;
      RECT 17.095 2.985 17.325 3.975 ;
      RECT 17.16 0.855 17.27 1.665 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.162 ;
  ANTENNAPARTIALMETALAREA 0.2528 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0706 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.84 1.82 1.845 2.1 ;
      RECT 1.305 1.67 1.84 2.14 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2188 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.945 2.38 1.18 2.66 ;
      RECT 0.605 2.21 0.945 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.22 -0.4 18.48 0.4 ;
      RECT 17.88 -0.4 18.22 1.485 ;
      RECT 16.78 -0.4 17.88 0.4 ;
      RECT 16.44 -0.4 16.78 1.485 ;
      RECT 15.34 -0.4 16.44 0.4 ;
      RECT 15 -0.4 15.34 0.95 ;
      RECT 14.04 -0.4 15 0.4 ;
      RECT 13.7 -0.4 14.04 1.55 ;
      RECT 11.44 -0.4 13.7 0.4 ;
      RECT 11.1 -0.4 11.44 0.575 ;
      RECT 9.45 -0.4 11.1 0.4 ;
      RECT 9.11 -0.4 9.45 1.32 ;
      RECT 6.89 -0.4 9.11 0.4 ;
      RECT 6.55 -0.4 6.89 1.32 ;
      RECT 3.97 -0.4 6.55 0.4 ;
      RECT 3.63 -0.4 3.97 1.28 ;
      RECT 1.25 -0.4 3.63 0.4 ;
      RECT 0.91 -0.4 1.25 0.575 ;
      RECT 0 -0.4 0.91 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.1 4.64 18.48 5.44 ;
      RECT 17.76 3.605 18.1 5.44 ;
      RECT 16.66 4.64 17.76 5.44 ;
      RECT 16.32 4.03 16.66 5.44 ;
      RECT 15.22 4.64 16.32 5.44 ;
      RECT 14.88 4.09 15.22 5.44 ;
      RECT 13.96 4.64 14.88 5.44 ;
      RECT 13.62 2.975 13.96 5.44 ;
      RECT 12.52 4.64 13.62 5.44 ;
      RECT 12.18 3.435 12.52 5.44 ;
      RECT 11.04 4.64 12.18 5.44 ;
      RECT 10.7 4.04 11.04 5.44 ;
      RECT 9.33 4.64 10.7 5.44 ;
      RECT 8.99 3.6 9.33 5.44 ;
      RECT 6.78 4.64 8.99 5.44 ;
      RECT 6.44 4.14 6.78 5.44 ;
      RECT 5.6 4.64 6.44 5.44 ;
      RECT 5.37 4.14 5.6 5.44 ;
      RECT 4.03 4.64 5.37 5.44 ;
      RECT 3.69 4.15 4.03 5.44 ;
      RECT 1.265 4.64 3.69 5.44 ;
      RECT 0.925 4.465 1.265 5.44 ;
      RECT 0 4.64 0.925 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 16.86 2.04 17.03 2.38 ;
      RECT 16.63 2.04 16.86 3.685 ;
      RECT 14.76 3.455 16.63 3.685 ;
      RECT 14.76 1.31 14.8 1.65 ;
      RECT 14.68 1.31 14.76 3.685 ;
      RECT 14.53 1.31 14.68 3.71 ;
      RECT 14.46 1.31 14.53 1.65 ;
      RECT 14.34 2.9 14.53 3.71 ;
      RECT 13.24 2.08 14.3 2.42 ;
      RECT 13.01 1.375 13.24 3.785 ;
      RECT 12.76 1.375 13.01 1.605 ;
      RECT 12.9 2.975 13.01 3.785 ;
      RECT 11.8 2.975 12.9 3.205 ;
      RECT 12.42 0.79 12.76 1.605 ;
      RECT 12.18 1.895 12.52 2.705 ;
      RECT 11.11 1.11 12.42 1.34 ;
      RECT 10.105 2.185 12.18 2.415 ;
      RECT 11.46 2.975 11.8 3.785 ;
      RECT 10.45 3.365 11.46 3.595 ;
      RECT 10.77 1 11.11 1.34 ;
      RECT 10.22 3.365 10.45 4.04 ;
      RECT 10.11 3.7 10.22 4.04 ;
      RECT 10.105 1.43 10.16 1.77 ;
      RECT 9.88 1.43 10.105 3.13 ;
      RECT 9.875 1.43 9.88 3.24 ;
      RECT 9.82 1.43 9.875 1.78 ;
      RECT 9.54 2.9 9.875 3.24 ;
      RECT 8.875 1.55 9.82 1.78 ;
      RECT 9.305 2.33 9.645 2.67 ;
      RECT 8.01 2.9 9.54 3.13 ;
      RECT 8.36 2.33 9.305 2.56 ;
      RECT 8.645 1.19 8.875 1.78 ;
      RECT 8.17 1.19 8.645 1.42 ;
      RECT 8.13 1.72 8.36 2.56 ;
      RECT 7.83 1.08 8.17 1.42 ;
      RECT 8.02 1.72 8.13 2.06 ;
      RECT 6.835 1.775 8.02 2.005 ;
      RECT 7.67 2.865 8.01 3.675 ;
      RECT 7.355 2.365 7.69 2.595 ;
      RECT 7.125 2.365 7.355 3.78 ;
      RECT 6.165 3.55 7.125 3.78 ;
      RECT 6.605 1.765 6.835 3.21 ;
      RECT 6.09 1.765 6.605 2.005 ;
      RECT 6.11 2.98 6.605 3.21 ;
      RECT 6.035 2.27 6.375 2.61 ;
      RECT 5.935 3.55 6.165 4.025 ;
      RECT 5.77 2.98 6.11 3.32 ;
      RECT 5.98 1.16 6.09 2.005 ;
      RECT 5.34 2.325 6.035 2.555 ;
      RECT 5.805 0.685 5.98 2.005 ;
      RECT 2.105 3.55 5.935 3.78 ;
      RECT 5.75 0.685 5.805 1.5 ;
      RECT 5.6 0.685 5.75 0.915 ;
      RECT 5.11 0.955 5.34 3.21 ;
      RECT 4.91 0.955 5.11 1.3 ;
      RECT 4.79 2.98 5.11 3.21 ;
      RECT 4.54 1.605 4.88 1.945 ;
      RECT 4.45 2.98 4.79 3.32 ;
      RECT 2.98 1.66 4.54 1.89 ;
      RECT 3.695 2.98 4.45 3.21 ;
      RECT 3.69 2.325 3.695 3.21 ;
      RECT 3.465 2.215 3.69 3.21 ;
      RECT 3.35 2.215 3.465 2.555 ;
      RECT 2.75 1.04 2.98 3.135 ;
      RECT 2.27 1.04 2.75 1.38 ;
      RECT 2.565 2.905 2.75 3.135 ;
      RECT 2.335 2.905 2.565 3.3 ;
      RECT 2.175 1.61 2.405 2.66 ;
      RECT 2.105 2.43 2.175 2.66 ;
      RECT 1.875 2.43 2.105 3.78 ;
      RECT 0.61 3.07 1.875 3.3 ;
      RECT 0.375 1.255 0.69 1.595 ;
      RECT 0.375 2.96 0.61 3.3 ;
      RECT 0.145 1.255 0.375 3.3 ;
  END
END DFFSX4

MACRO DFFSX2
  CLASS CORE ;
  FOREIGN DFFSX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.522 ;
  ANTENNAPARTIALMETALAREA 1.3956 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.4713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.085 4.005 9.685 4.355 ;
      RECT 3.93 4.005 9.085 4.235 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.0944 ;
  ANTENNAPARTIALMETALAREA 0.8972 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9909 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.86 1.26 12.325 1.54 ;
      RECT 11.63 0.63 11.86 2.94 ;
      RECT 11.37 0.63 11.63 0.97 ;
      RECT 11.58 2.635 11.63 2.94 ;
      RECT 11.36 2.635 11.58 3.05 ;
      RECT 11.24 2.71 11.36 3.05 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.44 ;
  ANTENNAPARTIALMETALAREA 1.3674 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.1251 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.415 1.325 13.645 3.115 ;
      RECT 13.34 1.26 13.415 3.115 ;
      RECT 13.23 1.26 13.34 1.555 ;
      RECT 13.02 2.885 13.34 3.115 ;
      RECT 12.89 0.745 13.23 1.555 ;
      RECT 12.68 2.885 13.02 4.165 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2034 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.29 2.36 1.805 2.755 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.2033 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9699 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.135 2.295 0.515 2.83 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.47 -0.4 13.86 0.4 ;
      RECT 12.13 -0.4 12.47 0.575 ;
      RECT 11.01 -0.4 12.13 0.4 ;
      RECT 10.67 -0.4 11.01 0.575 ;
      RECT 8.63 -0.4 10.67 0.4 ;
      RECT 8.29 -0.4 8.63 1.565 ;
      RECT 6.085 -0.4 8.29 0.4 ;
      RECT 5.855 -0.4 6.085 1.3 ;
      RECT 3.86 -0.4 5.855 0.4 ;
      RECT 3.52 -0.4 3.86 1.13 ;
      RECT 1.45 -0.4 3.52 0.4 ;
      RECT 1.11 -0.4 1.45 0.575 ;
      RECT 0 -0.4 1.11 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.3 4.64 13.86 5.44 ;
      RECT 11.96 3.865 12.3 5.44 ;
      RECT 10.33 4.64 11.96 5.44 ;
      RECT 9.99 3.445 10.33 5.44 ;
      RECT 9.98 3.445 9.99 3.785 ;
      RECT 8.84 4.64 9.99 5.44 ;
      RECT 8.5 4.465 8.84 5.44 ;
      RECT 6.36 4.64 8.5 5.44 ;
      RECT 6.02 4.465 6.36 5.44 ;
      RECT 5.1 4.64 6.02 5.44 ;
      RECT 4.76 4.465 5.1 5.44 ;
      RECT 3.7 4.64 4.76 5.44 ;
      RECT 3.36 4.465 3.7 5.44 ;
      RECT 1.31 4.64 3.36 5.44 ;
      RECT 0.97 4.465 1.31 5.44 ;
      RECT 0 4.64 0.97 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.45 2.07 12.67 2.41 ;
      RECT 12.22 2.07 12.45 3.545 ;
      RECT 11.04 3.315 12.22 3.545 ;
      RECT 11.01 1.345 11.17 1.685 ;
      RECT 11.01 3.315 11.04 3.78 ;
      RECT 10.78 1.345 11.01 3.78 ;
      RECT 10.7 3.44 10.78 3.78 ;
      RECT 10.405 2.015 10.515 2.355 ;
      RECT 10.175 1.795 10.405 3.125 ;
      RECT 9.91 1.795 10.175 2.025 ;
      RECT 9.6 2.895 10.175 3.125 ;
      RECT 9.57 1.335 9.91 2.025 ;
      RECT 9.5 2.255 9.84 2.665 ;
      RECT 9.26 2.895 9.6 3.705 ;
      RECT 8.33 1.795 9.57 2.025 ;
      RECT 7.68 2.435 9.5 2.665 ;
      RECT 7.99 1.795 8.33 2.205 ;
      RECT 7.625 2.435 7.68 3.775 ;
      RECT 7.395 1.405 7.625 3.775 ;
      RECT 7.305 1.405 7.395 1.75 ;
      RECT 7.34 3.545 7.395 3.775 ;
      RECT 7.11 2.54 7.145 2.88 ;
      RECT 6.88 2.54 7.11 3.775 ;
      RECT 6.645 1.735 7.06 2.075 ;
      RECT 2.82 3.545 6.88 3.775 ;
      RECT 6.415 1.53 6.645 3.03 ;
      RECT 5.625 1.53 6.415 1.76 ;
      RECT 5.86 2.8 6.415 3.03 ;
      RECT 5.165 1.99 6.17 2.33 ;
      RECT 5.52 2.8 5.86 3.14 ;
      RECT 5.395 0.84 5.625 1.76 ;
      RECT 5.22 0.84 5.395 1.07 ;
      RECT 4.88 0.635 5.22 1.07 ;
      RECT 4.935 1.44 5.165 3.315 ;
      RECT 3.55 3.085 4.935 3.315 ;
      RECT 4.09 0.635 4.88 0.865 ;
      RECT 4.54 2.445 4.65 2.785 ;
      RECT 4.31 2.125 4.54 2.785 ;
      RECT 2.83 2.125 4.31 2.355 ;
      RECT 3.32 2.59 3.55 3.315 ;
      RECT 3.21 2.59 3.32 2.93 ;
      RECT 2.825 0.815 2.83 3.115 ;
      RECT 2.6 0.76 2.825 3.115 ;
      RECT 2.48 3.545 2.82 4.06 ;
      RECT 2.485 0.76 2.6 1.1 ;
      RECT 2.54 2.885 2.6 3.115 ;
      RECT 2.2 2.885 2.54 3.225 ;
      RECT 0.98 3.545 2.48 3.775 ;
      RECT 2.03 1.725 2.37 2.065 ;
      RECT 0.98 1.78 2.03 2.01 ;
      RECT 0.75 1.78 0.98 3.775 ;
      RECT 0.525 1.78 0.75 2.01 ;
      RECT 0.55 3.45 0.75 3.775 ;
      RECT 0.21 3.45 0.55 3.79 ;
      RECT 0.295 1.19 0.525 2.01 ;
      RECT 0.185 1.19 0.295 1.53 ;
  END
END DFFSX2

MACRO DFFSX1
  CLASS CORE ;
  FOREIGN DFFSX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.54 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3348 ;
  ANTENNAPARTIALMETALAREA 0.2091 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9752 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.38 3.9 9.79 4.41 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6816 ;
  ANTENNAPARTIALMETALAREA 1.2856 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.8141 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.46 0.87 11.69 3.87 ;
      RECT 10.945 0.87 11.46 1.1 ;
      RECT 11.1 3.64 11.46 3.87 ;
      RECT 10.76 3.64 11.1 4.37 ;
      RECT 10.605 0.67 10.945 1.1 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.5605 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5811 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.325 2.63 12.36 3.21 ;
      RECT 12.095 1.25 12.325 3.21 ;
      RECT 11.96 1.25 12.095 1.59 ;
      RECT 12.02 2.63 12.095 3.21 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.205 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.435 1.08 1.845 1.58 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.3318 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.7172 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.955 2.965 1.105 3.195 ;
      RECT 0.725 2.575 0.955 3.195 ;
      RECT 0.555 2.575 0.725 2.805 ;
      RECT 0.215 2.465 0.555 2.805 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.685 -0.4 12.54 0.4 ;
      RECT 11.345 -0.4 11.685 0.575 ;
      RECT 10.22 -0.4 11.345 0.4 ;
      RECT 9.88 -0.4 10.22 0.96 ;
      RECT 8.56 -0.4 9.88 0.4 ;
      RECT 8.22 -0.4 8.56 0.575 ;
      RECT 6.165 -0.4 8.22 0.4 ;
      RECT 5.935 -0.4 6.165 1.01 ;
      RECT 4.04 -0.4 5.935 0.4 ;
      RECT 3.7 -0.4 4.04 1.11 ;
      RECT 1.545 -0.4 3.7 0.4 ;
      RECT 1.205 -0.4 1.545 0.575 ;
      RECT 0 -0.4 1.205 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.36 4.64 12.54 5.44 ;
      RECT 12.305 4.465 12.36 5.44 ;
      RECT 12.075 4.41 12.305 5.44 ;
      RECT 12.02 4.465 12.075 5.44 ;
      RECT 10.38 4.64 12.02 5.44 ;
      RECT 10.04 2.94 10.38 5.44 ;
      RECT 8.93 4.64 10.04 5.44 ;
      RECT 8.59 4.14 8.93 5.44 ;
      RECT 6.42 4.64 8.59 5.44 ;
      RECT 6.08 4.14 6.42 5.44 ;
      RECT 5.16 4.64 6.08 5.44 ;
      RECT 4.82 4.14 5.16 5.44 ;
      RECT 3.76 4.64 4.82 5.44 ;
      RECT 3.42 4.465 3.76 5.44 ;
      RECT 1.3 4.64 3.42 5.44 ;
      RECT 0.96 4.465 1.3 5.44 ;
      RECT 0 4.64 0.96 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 10.995 1.57 11.225 3.28 ;
      RECT 10.985 1.57 10.995 1.8 ;
      RECT 10.815 2.94 10.995 3.28 ;
      RECT 10.645 1.46 10.985 1.8 ;
      RECT 9.66 2.04 10.37 2.27 ;
      RECT 9.43 1.52 9.66 3.4 ;
      RECT 8.9 1.52 9.43 1.75 ;
      RECT 9.32 3.06 9.43 3.4 ;
      RECT 7.74 2.465 9.2 2.695 ;
      RECT 8.56 1.405 8.9 1.75 ;
      RECT 8.22 1.405 8.56 1.645 ;
      RECT 7.88 1.305 8.22 1.645 ;
      RECT 7.63 2.465 7.74 3.65 ;
      RECT 7.4 1.54 7.63 3.65 ;
      RECT 7.325 1.54 7.4 1.77 ;
      RECT 7.165 4.02 7.37 4.36 ;
      RECT 7.095 1.43 7.325 1.77 ;
      RECT 6.935 3.67 7.165 4.36 ;
      RECT 6.84 2.335 7.1 2.675 ;
      RECT 2.88 3.67 6.935 3.9 ;
      RECT 6.61 1.24 6.84 3.31 ;
      RECT 5.705 1.24 6.61 1.47 ;
      RECT 5.865 3.08 6.61 3.31 ;
      RECT 5.245 2.165 6.375 2.505 ;
      RECT 5.635 3.08 5.865 3.42 ;
      RECT 5.475 0.78 5.705 1.47 ;
      RECT 5.385 0.78 5.475 1.01 ;
      RECT 5.38 0.675 5.385 1.01 ;
      RECT 5.04 0.67 5.38 1.01 ;
      RECT 5.015 1.42 5.245 3.23 ;
      RECT 4.27 0.675 5.04 0.905 ;
      RECT 4.56 3 5.015 3.23 ;
      RECT 4.725 2.395 4.73 2.735 ;
      RECT 4.39 2.18 4.725 2.735 ;
      RECT 4.22 3 4.56 3.34 ;
      RECT 2.91 2.18 4.39 2.41 ;
      RECT 3.6 3 4.22 3.23 ;
      RECT 3.37 2.64 3.6 3.23 ;
      RECT 3.26 2.64 3.37 2.98 ;
      RECT 2.68 0.74 2.91 3.115 ;
      RECT 2.54 3.56 2.88 4.14 ;
      RECT 2.565 0.74 2.68 1.08 ;
      RECT 2.6 2.885 2.68 3.115 ;
      RECT 2.26 2.885 2.6 3.225 ;
      RECT 1.905 3.56 2.54 3.79 ;
      RECT 2.105 1.82 2.445 2.16 ;
      RECT 1.905 1.93 2.105 2.16 ;
      RECT 1.655 1.93 1.905 3.79 ;
      RECT 0.53 1.93 1.655 2.16 ;
      RECT 0.195 3.45 1.655 3.79 ;
      RECT 0.3 1.19 0.53 2.16 ;
      RECT 0.19 1.19 0.3 1.53 ;
  END
END DFFSX1

MACRO DFFRHQXL
  CLASS CORE ;
  FOREIGN DFFRHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2765 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.61 2.91 12.4 3.26 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6804 ;
  ANTENNAPARTIALMETALAREA 0.9661 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5633 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.645 3.715 13.66 4.055 ;
      RECT 13.415 1.305 13.645 4.055 ;
      RECT 12.755 1.305 13.415 1.535 ;
      RECT 13.32 3.715 13.415 4.055 ;
      RECT 12.65 1.26 12.755 1.535 ;
      RECT 12.31 1.195 12.65 1.535 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2064 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.36 1.68 1.84 2.11 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9964 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.63 2.17 1.105 2.635 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.87 -0.4 13.86 0.4 ;
      RECT 12.53 -0.4 12.87 0.575 ;
      RECT 11.365 -0.4 12.53 0.4 ;
      RECT 11.025 -0.4 11.365 0.575 ;
      RECT 9.765 -0.4 11.025 0.4 ;
      RECT 9.425 -0.4 9.765 0.575 ;
      RECT 6.79 -0.4 9.425 0.4 ;
      RECT 6.45 -0.4 6.79 1.16 ;
      RECT 4.1 -0.4 6.45 0.4 ;
      RECT 5.4 1.47 5.51 1.81 ;
      RECT 5.17 1.205 5.4 1.81 ;
      RECT 4.1 1.205 5.17 1.435 ;
      RECT 3.76 -0.4 4.1 1.435 ;
      RECT 1.48 -0.4 3.76 0.4 ;
      RECT 1.14 -0.4 1.48 0.575 ;
      RECT 0 -0.4 1.14 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.38 4.64 13.86 5.44 ;
      RECT 12.04 3.49 12.38 5.44 ;
      RECT 11.28 3.49 12.04 3.72 ;
      RECT 10.09 4.64 12.04 5.44 ;
      RECT 11.05 3.205 11.28 3.72 ;
      RECT 10.94 3.205 11.05 3.545 ;
      RECT 9.675 4.465 10.09 5.44 ;
      RECT 7.135 4.64 9.675 5.44 ;
      RECT 6.795 4.465 7.135 5.44 ;
      RECT 4.04 4.64 6.795 5.44 ;
      RECT 3.7 4 4.04 5.44 ;
      RECT 1.48 4.64 3.7 5.44 ;
      RECT 1.14 3.885 1.48 5.44 ;
      RECT 0 4.64 1.14 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 11.8 1.78 13.18 2.01 ;
      RECT 11.245 2.45 12.69 2.68 ;
      RECT 11.57 0.855 11.8 2.01 ;
      RECT 11.24 3.98 11.58 4.32 ;
      RECT 10.125 0.855 11.57 1.085 ;
      RECT 10.905 1.315 11.245 2.68 ;
      RECT 10.625 3.98 11.24 4.21 ;
      RECT 10.625 2.21 10.905 2.68 ;
      RECT 10.585 2.21 10.625 4.21 ;
      RECT 10.395 2.405 10.585 4.21 ;
      RECT 9.96 1.465 10.44 1.695 ;
      RECT 5.785 3.945 10.395 4.175 ;
      RECT 9.755 0.855 10.125 1.235 ;
      RECT 9.73 1.465 9.96 3.55 ;
      RECT 9.225 1.005 9.755 1.235 ;
      RECT 9.62 2.58 9.73 3.55 ;
      RECT 9.455 2.58 9.62 2.93 ;
      RECT 8.995 1.005 9.225 3.6 ;
      RECT 8.4 1.005 8.995 1.255 ;
      RECT 8.67 3.37 8.995 3.6 ;
      RECT 8.48 1.61 8.715 1.95 ;
      RECT 8.33 3.37 8.67 3.71 ;
      RECT 8.25 1.61 8.48 3.055 ;
      RECT 8.06 1.005 8.4 1.365 ;
      RECT 7.795 1.595 8.02 3.71 ;
      RECT 7.79 1.01 7.795 3.71 ;
      RECT 7.565 1.01 7.79 1.825 ;
      RECT 7.61 3.37 7.79 3.71 ;
      RECT 7.26 1.01 7.565 1.35 ;
      RECT 7.335 2.28 7.56 2.62 ;
      RECT 7.105 1.63 7.335 3.58 ;
      RECT 6.34 1.63 7.105 1.86 ;
      RECT 6.63 3.35 7.105 3.58 ;
      RECT 6.635 2.175 6.865 2.915 ;
      RECT 4.815 2.175 6.635 2.405 ;
      RECT 6.29 3.35 6.63 3.69 ;
      RECT 6.205 1.52 6.34 1.86 ;
      RECT 5.975 0.685 6.205 1.86 ;
      RECT 4.7 0.685 5.975 0.915 ;
      RECT 5.555 2.635 5.785 4.175 ;
      RECT 5.325 2.635 5.555 2.975 ;
      RECT 4.585 1.67 4.815 3.68 ;
      RECT 4.36 0.63 4.7 0.97 ;
      RECT 4.37 1.67 4.585 2.01 ;
      RECT 4.41 3.34 4.585 3.68 ;
      RECT 3.695 1.78 4.37 2.01 ;
      RECT 4.12 2.58 4.35 2.945 ;
      RECT 2.935 2.715 4.12 2.945 ;
      RECT 3.465 1.78 3.695 2.37 ;
      RECT 3.355 2.03 3.465 2.37 ;
      RECT 2.83 3.74 3.17 4.08 ;
      RECT 2.76 1.24 2.935 2.945 ;
      RECT 2.3 3.74 2.83 3.97 ;
      RECT 2.705 1.24 2.76 3.325 ;
      RECT 2.7 1.24 2.705 1.47 ;
      RECT 2.53 2.715 2.705 3.325 ;
      RECT 2.36 1.13 2.7 1.47 ;
      RECT 2.3 1.81 2.465 2.15 ;
      RECT 2.07 1.81 2.3 3.97 ;
      RECT 0.83 3 2.07 3.23 ;
      RECT 0.49 2.89 0.83 3.23 ;
      RECT 0.4 1.34 0.625 1.71 ;
      RECT 0.4 2.89 0.49 3.12 ;
      RECT 0.17 1.34 0.4 3.12 ;
  END
END DFFRHQXL

MACRO DFFRHQX4
  CLASS CORE ;
  FOREIGN DFFRHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 21.12 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRHQXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.738 ;
  ANTENNAPARTIALMETALAREA 0.25 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.485 1.82 14.965 2.1 ;
      RECT 14.145 1.78 14.485 2.12 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.6352 ;
  ANTENNAPARTIALMETALAREA 2.6363 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.9799 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.525 2.965 20.865 3.835 ;
      RECT 20.32 2.965 20.525 3.22 ;
      RECT 19.94 1.415 20.32 3.22 ;
      RECT 19.5 1.415 19.94 1.645 ;
      RECT 18.305 2.99 19.94 3.22 ;
      RECT 19.16 0.785 19.5 1.645 ;
      RECT 18.06 1.415 19.16 1.645 ;
      RECT 17.965 2.99 18.305 3.835 ;
      RECT 17.72 0.785 18.06 1.645 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3348 ;
  ANTENNAPARTIALMETALAREA 0.2577 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3303 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.24 2.075 1.47 2.66 ;
      RECT 0.8 2.38 1.24 2.66 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.4932 ;
  ANTENNAPARTIALMETALAREA 0.2288 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.785 0.855 2.105 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.26 -0.4 21.12 0.4 ;
      RECT 19.92 -0.4 20.26 1.1 ;
      RECT 18.78 -0.4 19.92 0.4 ;
      RECT 18.44 -0.4 18.78 1.185 ;
      RECT 17.325 -0.4 18.44 0.4 ;
      RECT 16.985 -0.4 17.325 1.565 ;
      RECT 15.485 -0.4 16.985 0.4 ;
      RECT 15.145 -0.4 15.485 0.575 ;
      RECT 14.005 -0.4 15.145 0.4 ;
      RECT 13.665 -0.4 14.005 1.32 ;
      RECT 8.465 -0.4 13.665 0.4 ;
      RECT 8.125 -0.4 8.465 1.32 ;
      RECT 7.025 -0.4 8.125 0.4 ;
      RECT 6.685 -0.4 7.025 1.49 ;
      RECT 5.365 -0.4 6.685 0.4 ;
      RECT 5.365 1.26 5.405 1.6 ;
      RECT 5.065 -0.4 5.365 1.6 ;
      RECT 3.925 -0.4 5.065 0.4 ;
      RECT 3.585 -0.4 3.925 0.97 ;
      RECT 1.31 -0.4 3.585 0.4 ;
      RECT 0.97 -0.4 1.31 0.575 ;
      RECT 0 -0.4 0.97 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.585 4.64 21.12 5.44 ;
      RECT 19.245 3.45 19.585 5.44 ;
      RECT 16.97 4.64 19.245 5.44 ;
      RECT 16.74 3.11 16.97 5.44 ;
      RECT 15.325 4.64 16.74 5.44 ;
      RECT 14.985 4.465 15.325 5.44 ;
      RECT 13.625 4.64 14.985 5.44 ;
      RECT 13.395 4.08 13.625 5.44 ;
      RECT 8.685 4.64 13.395 5.44 ;
      RECT 8.345 4.465 8.685 5.44 ;
      RECT 7.16 4.64 8.345 5.44 ;
      RECT 6.93 4.04 7.16 5.44 ;
      RECT 5.735 4.64 6.93 5.44 ;
      RECT 5.395 4.465 5.735 5.44 ;
      RECT 3.845 4.64 5.395 5.44 ;
      RECT 3.505 4.465 3.845 5.44 ;
      RECT 1.2 4.64 3.505 5.44 ;
      RECT 1.2 3.485 1.255 3.825 ;
      RECT 0.97 3.485 1.2 5.44 ;
      RECT 0.915 3.485 0.97 3.825 ;
      RECT 0 4.64 0.97 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 18.88 2.045 19.22 2.385 ;
      RECT 16.785 2.125 18.88 2.355 ;
      RECT 16.755 2.125 16.785 2.55 ;
      RECT 16.525 0.805 16.755 2.55 ;
      RECT 14.725 0.805 16.525 1.035 ;
      RECT 16.51 2.125 16.525 2.55 ;
      RECT 16.28 2.125 16.51 4.14 ;
      RECT 16.065 1.265 16.295 1.605 ;
      RECT 14.49 3.91 16.28 4.14 ;
      RECT 15.565 1.375 16.065 1.605 ;
      RECT 15.82 2.2 16.05 3.57 ;
      RECT 14.66 3.34 15.82 3.57 ;
      RECT 15.335 1.375 15.565 3.11 ;
      RECT 13.745 2.36 15.335 2.59 ;
      RECT 14.385 0.805 14.725 1.33 ;
      RECT 14.43 3.16 14.66 3.57 ;
      RECT 14.15 3.91 14.49 4.25 ;
      RECT 13.135 3.16 14.43 3.39 ;
      RECT 13.92 3.62 14.15 4.14 ;
      RECT 13.16 3.62 13.92 3.85 ;
      RECT 13.515 2.245 13.745 2.59 ;
      RECT 13.265 2.245 13.515 2.475 ;
      RECT 12.925 2.135 13.265 2.475 ;
      RECT 12.93 3.62 13.16 4.365 ;
      RECT 12.905 2.78 13.135 3.39 ;
      RECT 9.145 4.135 12.93 4.365 ;
      RECT 12.51 2.78 12.905 3.01 ;
      RECT 12.615 3.28 12.67 3.62 ;
      RECT 12.51 1.1 12.645 1.44 ;
      RECT 12.33 3.28 12.615 3.845 ;
      RECT 12.28 0.675 12.51 3.01 ;
      RECT 9.725 3.615 12.33 3.845 ;
      RECT 11.205 0.675 12.28 0.905 ;
      RECT 12.055 2.635 12.28 3.01 ;
      RECT 10.82 2.635 12.055 2.865 ;
      RECT 11.815 1.14 11.925 1.48 ;
      RECT 11.585 1.14 11.815 1.84 ;
      RECT 10.485 1.61 11.585 1.84 ;
      RECT 10.185 3.095 11.58 3.325 ;
      RECT 10.865 0.675 11.205 1.38 ;
      RECT 9.385 0.675 10.865 0.905 ;
      RECT 10.535 2.52 10.82 2.865 ;
      RECT 10.48 2.52 10.535 2.86 ;
      RECT 10.145 1.14 10.485 1.84 ;
      RECT 10.12 2.905 10.185 3.325 ;
      RECT 10.12 1.31 10.145 1.84 ;
      RECT 9.955 1.31 10.12 3.325 ;
      RECT 9.89 1.31 9.955 3.19 ;
      RECT 9.185 1.31 9.89 1.54 ;
      RECT 9.715 2.85 9.89 3.19 ;
      RECT 9.495 3.425 9.725 3.845 ;
      RECT 8.65 2.905 9.715 3.135 ;
      RECT 9.43 1.77 9.66 2.435 ;
      RECT 8.08 3.425 9.495 3.655 ;
      RECT 8.08 2.205 9.43 2.435 ;
      RECT 8.845 1.31 9.185 1.785 ;
      RECT 8.915 4.005 9.145 4.365 ;
      RECT 7.62 4.005 8.915 4.235 ;
      RECT 7.745 1.555 8.845 1.785 ;
      RECT 8.31 2.77 8.65 3.135 ;
      RECT 7.85 2.205 8.08 3.655 ;
      RECT 7.15 2.205 7.85 2.435 ;
      RECT 7.515 1.15 7.745 1.785 ;
      RECT 7.39 3.295 7.62 4.235 ;
      RECT 7.405 1.15 7.515 1.49 ;
      RECT 6.535 3.295 7.39 3.525 ;
      RECT 7.095 2.205 7.15 3.06 ;
      RECT 6.865 1.775 7.095 3.06 ;
      RECT 6.3 1.775 6.865 2.005 ;
      RECT 6.81 2.72 6.865 3.06 ;
      RECT 6.4 3.88 6.63 4.225 ;
      RECT 6.305 2.235 6.535 3.525 ;
      RECT 3.04 3.995 6.4 4.225 ;
      RECT 5.335 2.235 6.305 2.465 ;
      RECT 6.19 1.26 6.3 2.005 ;
      RECT 5.96 0.675 6.19 2.005 ;
      RECT 5.735 2.93 6.075 3.3 ;
      RECT 5.595 0.675 5.96 0.905 ;
      RECT 4.765 2.93 5.735 3.16 ;
      RECT 4.995 2.11 5.335 2.465 ;
      RECT 4.535 1.14 4.765 3.16 ;
      RECT 4.345 1.14 4.535 1.48 ;
      RECT 4.38 2.93 4.535 3.16 ;
      RECT 4.04 2.93 4.38 3.27 ;
      RECT 3.945 2.04 4.285 2.64 ;
      RECT 3.615 2.93 4.04 3.16 ;
      RECT 2.735 2.04 3.945 2.27 ;
      RECT 3.275 2.57 3.615 3.16 ;
      RECT 2.81 2.67 3.04 4.225 ;
      RECT 2.645 2.67 2.81 3.065 ;
      RECT 1.95 3.995 2.81 4.225 ;
      RECT 2.505 0.9 2.735 2.27 ;
      RECT 2.415 3.42 2.55 3.76 ;
      RECT 2.305 0.9 2.505 1.24 ;
      RECT 2.415 2.04 2.505 2.27 ;
      RECT 2.185 2.04 2.415 3.76 ;
      RECT 1.95 1.47 2.275 1.81 ;
      RECT 1.72 1.275 1.95 4.225 ;
      RECT 0.535 1.275 1.72 1.505 ;
      RECT 0.535 2.89 1.72 3.245 ;
      RECT 0.195 0.695 0.535 1.505 ;
      RECT 0.195 2.89 0.535 4.17 ;
  END
END DFFRHQX4

MACRO DFFRHQX2
  CLASS CORE ;
  FOREIGN DFFRHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRHQXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.414 ;
  ANTENNAPARTIALMETALAREA 0.2942 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1501 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.415 2.655 13.95 3.205 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.296 ;
  ANTENNAPARTIALMETALAREA 1.4696 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.254 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.16 1.21 16.39 3.105 ;
      RECT 15.03 1.21 16.16 1.44 ;
      RECT 15.7 2.875 16.16 3.105 ;
      RECT 15.36 2.875 15.7 4.03 ;
      RECT 14.69 0.635 15.03 1.445 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.198 ;
  ANTENNAPARTIALMETALAREA 0.2354 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0706 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.645 1.72 1.84 2.085 ;
      RECT 1.28 1.72 1.645 2.14 ;
      RECT 1.25 1.72 1.28 2.085 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.306 ;
  ANTENNAPARTIALMETALAREA 0.2107 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0123 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.02 2.38 1.105 2.635 ;
      RECT 0.6 2.23 1.02 2.68 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.79 -0.4 17.16 0.4 ;
      RECT 15.45 -0.4 15.79 0.575 ;
      RECT 14.045 -0.4 15.45 0.4 ;
      RECT 13.105 -0.4 14.045 0.575 ;
      RECT 11.76 -0.4 13.105 0.4 ;
      RECT 11.42 -0.4 11.76 0.575 ;
      RECT 7.845 -0.4 11.42 0.4 ;
      RECT 7.505 -0.4 7.845 1.29 ;
      RECT 3.95 -0.4 7.505 0.4 ;
      RECT 5.34 1.435 5.45 1.775 ;
      RECT 5.11 1.205 5.34 1.775 ;
      RECT 3.95 1.205 5.11 1.435 ;
      RECT 3.61 -0.4 3.95 1.435 ;
      RECT 1.325 -0.4 3.61 0.4 ;
      RECT 0.985 -0.4 1.325 0.575 ;
      RECT 0 -0.4 0.985 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.98 4.64 17.16 5.44 ;
      RECT 16.64 3.295 16.98 5.44 ;
      RECT 14.33 4.64 16.64 5.44 ;
      RECT 13.99 4.465 14.33 5.44 ;
      RECT 12.93 4.64 13.99 5.44 ;
      RECT 12.59 4.465 12.93 5.44 ;
      RECT 11.745 4.64 12.59 5.44 ;
      RECT 11.305 4.465 11.745 5.44 ;
      RECT 7.865 4.64 11.305 5.44 ;
      RECT 7.525 4.465 7.865 5.44 ;
      RECT 4.04 4.64 7.525 5.44 ;
      RECT 3.7 4 4.04 5.44 ;
      RECT 1.54 4.64 3.7 5.44 ;
      RECT 1.2 3.835 1.54 5.44 ;
      RECT 0 4.64 1.2 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.35 2.305 15.93 2.645 ;
      RECT 15.12 1.675 15.35 2.645 ;
      RECT 14.155 1.675 15.12 1.905 ;
      RECT 14.39 2.17 14.73 2.57 ;
      RECT 13.69 2.17 14.39 2.4 ;
      RECT 13.925 0.865 14.155 1.905 ;
      RECT 12.305 0.865 13.925 1.095 ;
      RECT 13.45 3.61 13.79 3.95 ;
      RECT 13.35 1.48 13.69 2.4 ;
      RECT 12.95 3.61 13.45 3.84 ;
      RECT 12.95 2.17 13.35 2.4 ;
      RECT 12.84 2.17 12.95 3.84 ;
      RECT 12.61 2.17 12.84 4.175 ;
      RECT 12.29 1.41 12.63 1.75 ;
      RECT 10.425 3.945 12.61 4.175 ;
      RECT 11.95 0.865 12.305 1.145 ;
      RECT 11.91 1.52 12.29 1.75 ;
      RECT 10.395 0.865 11.95 1.095 ;
      RECT 11.57 1.52 11.91 3.5 ;
      RECT 11.565 1.52 11.57 2.88 ;
      RECT 11.29 2.54 11.565 2.88 ;
      RECT 10.57 1.51 10.68 1.85 ;
      RECT 10.34 1.51 10.57 3 ;
      RECT 10.195 3.945 10.425 4.365 ;
      RECT 10.055 0.66 10.395 1.095 ;
      RECT 10.19 2.66 10.34 3 ;
      RECT 8.325 4.135 10.195 4.365 ;
      RECT 9.965 3.34 10.16 3.68 ;
      RECT 9.29 0.865 10.055 1.095 ;
      RECT 9.96 1.42 10.015 1.76 ;
      RECT 9.96 3.34 9.965 3.845 ;
      RECT 9.73 1.42 9.96 3.845 ;
      RECT 9.675 1.42 9.73 1.76 ;
      RECT 8.785 3.615 9.73 3.845 ;
      RECT 9.29 2.96 9.44 3.3 ;
      RECT 9.06 0.865 9.29 3.3 ;
      RECT 8.95 1.42 9.06 1.76 ;
      RECT 8.66 3.365 8.785 3.845 ;
      RECT 8.565 1.52 8.66 3.845 ;
      RECT 8.555 1.21 8.565 3.845 ;
      RECT 8.43 1.21 8.555 3.71 ;
      RECT 8.225 1.21 8.43 1.75 ;
      RECT 8.38 3.37 8.43 3.71 ;
      RECT 7.34 3.425 8.38 3.655 ;
      RECT 8.095 3.945 8.325 4.365 ;
      RECT 7.07 1.52 8.225 1.75 ;
      RECT 7.97 1.98 8.2 3.135 ;
      RECT 5.66 3.945 8.095 4.175 ;
      RECT 6.605 1.98 7.97 2.21 ;
      RECT 6.64 2.905 7.97 3.135 ;
      RECT 6.145 2.445 7.58 2.675 ;
      RECT 7 3.37 7.34 3.71 ;
      RECT 6.84 1.06 7.07 1.75 ;
      RECT 6.41 2.905 6.64 3.545 ;
      RECT 6.375 1.33 6.605 2.21 ;
      RECT 6.3 3.205 6.41 3.545 ;
      RECT 6.255 1.33 6.375 1.56 ;
      RECT 6.145 1.22 6.255 1.56 ;
      RECT 5.915 0.74 6.145 1.56 ;
      RECT 5.915 2.005 6.145 2.675 ;
      RECT 4.6 0.74 5.915 0.97 ;
      RECT 4.795 2.005 5.915 2.235 ;
      RECT 5.66 2.55 5.665 2.89 ;
      RECT 5.43 2.55 5.66 4.175 ;
      RECT 5.325 2.55 5.43 2.89 ;
      RECT 4.65 1.78 4.795 3.68 ;
      RECT 4.565 1.67 4.65 3.68 ;
      RECT 4.26 0.63 4.6 0.97 ;
      RECT 4.31 1.67 4.565 2.01 ;
      RECT 4.415 3.34 4.565 3.68 ;
      RECT 3.995 2.55 4.335 2.945 ;
      RECT 3.665 1.78 4.31 2.01 ;
      RECT 2.895 2.715 3.995 2.945 ;
      RECT 3.435 1.78 3.665 2.48 ;
      RECT 3.325 2.14 3.435 2.48 ;
      RECT 3.05 3.79 3.105 4.13 ;
      RECT 2.765 3.785 3.05 4.13 ;
      RECT 2.665 1.395 2.895 3.325 ;
      RECT 2.305 3.785 2.765 4.015 ;
      RECT 2.585 1.395 2.665 1.625 ;
      RECT 2.535 2.93 2.665 3.325 ;
      RECT 2.245 0.815 2.585 1.625 ;
      RECT 2.075 1.855 2.305 4.015 ;
      RECT 0.78 2.91 2.075 3.14 ;
      RECT 0.44 2.91 0.78 3.72 ;
      RECT 0.36 1.195 0.665 1.535 ;
      RECT 0.36 2.91 0.44 3.14 ;
      RECT 0.13 1.195 0.36 3.14 ;
  END
END DFFRHQX2

MACRO DFFRHQX1
  CLASS CORE ;
  FOREIGN DFFRHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRHQXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2628 ;
  ANTENNAPARTIALMETALAREA 0.2765 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.61 2.91 12.4 3.26 ;
     END
  END RN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.924 ;
  ANTENNAPARTIALMETALAREA 1.2268 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.406 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.63 1.245 13.645 3.195 ;
      RECT 13.415 1.245 13.63 4.29 ;
      RECT 12.57 1.245 13.415 1.475 ;
      RECT 13.34 2.965 13.415 4.29 ;
      RECT 13.29 3.48 13.34 4.29 ;
      RECT 12.34 0.73 12.57 1.475 ;
      RECT 12.23 0.73 12.34 1.07 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2708 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4363 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.615 1.285 1.765 1.515 ;
      RECT 1.615 1.81 1.62 2.15 ;
      RECT 1.385 1.285 1.615 2.15 ;
      RECT 1.28 1.81 1.385 2.15 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.216 ;
  ANTENNAPARTIALMETALAREA 0.2091 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.9 2.405 1.105 2.66 ;
      RECT 0.58 2.17 0.9 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.29 -0.4 13.86 0.4 ;
      RECT 12.95 -0.4 13.29 0.95 ;
      RECT 11.805 -0.4 12.95 0.4 ;
      RECT 10.865 -0.4 11.805 0.575 ;
      RECT 9.725 -0.4 10.865 0.4 ;
      RECT 9.385 -0.4 9.725 0.575 ;
      RECT 6.795 -0.4 9.385 0.4 ;
      RECT 6.455 -0.4 6.795 1.13 ;
      RECT 4.02 -0.4 6.455 0.4 ;
      RECT 5.36 1.48 5.47 1.82 ;
      RECT 5.13 1.205 5.36 1.82 ;
      RECT 4.02 1.205 5.13 1.435 ;
      RECT 3.68 -0.4 4.02 1.435 ;
      RECT 1.295 -0.4 3.68 0.4 ;
      RECT 0.955 -0.4 1.295 1.045 ;
      RECT 0 -0.4 0.955 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.35 4.64 13.86 5.44 ;
      RECT 12.01 3.52 12.35 5.44 ;
      RECT 11.28 3.535 12.01 3.765 ;
      RECT 10.09 4.64 12.01 5.44 ;
      RECT 11.05 2.93 11.28 3.765 ;
      RECT 10.94 2.93 11.05 3.27 ;
      RECT 9.675 4.465 10.09 5.44 ;
      RECT 7.215 4.64 9.675 5.44 ;
      RECT 6.8 4.465 7.215 5.44 ;
      RECT 4.04 4.64 6.8 5.44 ;
      RECT 3.7 3.98 4.04 5.44 ;
      RECT 1.58 4.64 3.7 5.44 ;
      RECT 1.24 3.8 1.58 5.44 ;
      RECT 0 4.64 1.24 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.81 1.71 13.15 2.05 ;
      RECT 11.76 1.71 12.81 1.94 ;
      RECT 11.24 2.45 12.69 2.68 ;
      RECT 11.53 0.865 11.76 1.94 ;
      RECT 11.285 4 11.625 4.34 ;
      RECT 10.085 0.865 11.53 1.095 ;
      RECT 10.705 4 11.285 4.23 ;
      RECT 10.925 1.375 11.24 2.68 ;
      RECT 10.865 1.375 10.925 1.715 ;
      RECT 10.705 2.21 10.925 2.68 ;
      RECT 10.585 2.21 10.705 4.23 ;
      RECT 10.475 2.405 10.585 4.23 ;
      RECT 10.47 3.945 10.475 4.23 ;
      RECT 5.785 3.945 10.47 4.175 ;
      RECT 10.06 1.41 10.4 1.75 ;
      RECT 9.715 0.865 10.085 1.145 ;
      RECT 10.04 1.52 10.06 1.75 ;
      RECT 9.81 1.52 10.04 3.5 ;
      RECT 9.62 2.58 9.81 3.5 ;
      RECT 9.225 0.865 9.715 1.095 ;
      RECT 9.455 2.58 9.62 2.93 ;
      RECT 8.995 0.865 9.225 3.6 ;
      RECT 8.305 0.865 8.995 1.105 ;
      RECT 8.67 3.37 8.995 3.6 ;
      RECT 8.48 1.605 8.675 1.945 ;
      RECT 8.33 3.37 8.67 3.71 ;
      RECT 8.335 1.605 8.48 3.055 ;
      RECT 8.25 1.61 8.335 3.055 ;
      RECT 8.075 0.865 8.305 1.275 ;
      RECT 7.95 1.595 8.02 3.705 ;
      RECT 7.815 1.595 7.95 3.71 ;
      RECT 7.79 1.12 7.815 3.71 ;
      RECT 7.585 1.12 7.79 1.825 ;
      RECT 7.61 3.37 7.79 3.71 ;
      RECT 7.56 1.12 7.585 1.35 ;
      RECT 7.22 1.01 7.56 1.35 ;
      RECT 7.335 2.3 7.56 2.705 ;
      RECT 7.105 1.64 7.335 3.58 ;
      RECT 6.3 1.64 7.105 1.87 ;
      RECT 6.63 3.35 7.105 3.58 ;
      RECT 6.635 2.175 6.865 2.915 ;
      RECT 4.865 2.175 6.635 2.405 ;
      RECT 6.29 3.35 6.63 3.69 ;
      RECT 6.165 1.53 6.3 1.87 ;
      RECT 5.935 0.74 6.165 1.87 ;
      RECT 4.66 0.74 5.935 0.97 ;
      RECT 5.555 2.635 5.785 4.175 ;
      RECT 5.32 2.635 5.555 2.975 ;
      RECT 4.67 1.78 4.865 3.68 ;
      RECT 4.635 1.67 4.67 3.68 ;
      RECT 4.32 0.63 4.66 0.97 ;
      RECT 4.33 1.67 4.635 2.01 ;
      RECT 4.41 3.34 4.635 3.68 ;
      RECT 4.065 2.58 4.405 2.945 ;
      RECT 3.63 1.78 4.33 2.01 ;
      RECT 2.895 2.715 4.065 2.945 ;
      RECT 3.4 1.78 3.63 2.37 ;
      RECT 3.29 2.03 3.4 2.37 ;
      RECT 2.83 3.74 3.17 4.08 ;
      RECT 2.85 1.045 2.895 2.945 ;
      RECT 2.665 1.045 2.85 3.325 ;
      RECT 2.28 3.74 2.83 3.97 ;
      RECT 2.66 1.045 2.665 1.275 ;
      RECT 2.615 2.715 2.665 3.325 ;
      RECT 2.32 0.935 2.66 1.275 ;
      RECT 2.51 2.985 2.615 3.325 ;
      RECT 2.28 1.83 2.335 2.17 ;
      RECT 2.05 1.83 2.28 3.97 ;
      RECT 1.995 1.83 2.05 2.17 ;
      RECT 0.78 2.89 2.05 3.12 ;
      RECT 0.44 2.89 0.78 3.23 ;
      RECT 0.35 1.28 0.52 1.62 ;
      RECT 0.35 2.89 0.44 3.12 ;
      RECT 0.12 1.28 0.35 3.12 ;
  END
END DFFRHQX1

MACRO DFFRXL
  CLASS CORE ;
  FOREIGN DFFRXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.18 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2142 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.97 2.86 4.48 3.28 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5343 ;
  ANTENNAPARTIALMETALAREA 1.393 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.2434 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.01 0.865 14.24 3.755 ;
      RECT 13.41 0.865 14.01 1.095 ;
      RECT 13.695 3.525 14.01 3.755 ;
      RECT 13.645 3.525 13.695 4.035 ;
      RECT 13.315 3.5 13.645 4.035 ;
      RECT 13.07 0.635 13.41 1.095 ;
      RECT 13.25 3.805 13.315 4.035 ;
      RECT 12.91 3.805 13.25 4.23 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 0.8116 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5722 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.835 1.82 15.04 2.1 ;
      RECT 14.835 3.62 14.92 3.96 ;
      RECT 14.82 1.82 14.835 3.96 ;
      RECT 14.605 1.265 14.82 3.96 ;
      RECT 14.475 1.265 14.605 2.075 ;
      RECT 14.58 3.62 14.605 3.96 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2122 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0653 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.74 1.96 2.08 ;
      RECT 1.62 1.74 1.765 2.105 ;
      RECT 1.32 1.795 1.62 2.105 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3115 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2031 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.55 1.265 3.22 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.14 -0.4 15.18 0.4 ;
      RECT 13.8 -0.4 14.14 0.575 ;
      RECT 12.53 -0.4 13.8 0.4 ;
      RECT 12.19 -0.4 12.53 0.95 ;
      RECT 10.77 -0.4 12.19 0.4 ;
      RECT 10.43 -0.4 10.77 1.3 ;
      RECT 6.17 -0.4 10.43 0.4 ;
      RECT 7.87 1.42 7.88 1.76 ;
      RECT 7.54 1.205 7.87 1.76 ;
      RECT 6.58 1.205 7.54 1.435 ;
      RECT 6.24 1.205 6.58 1.56 ;
      RECT 6.17 1.205 6.24 1.505 ;
      RECT 5.94 -0.4 6.17 1.505 ;
      RECT 4.655 -0.4 5.94 0.4 ;
      RECT 4.315 -0.4 4.655 0.96 ;
      RECT 1.555 -0.4 4.315 0.4 ;
      RECT 1.215 -0.4 1.555 0.575 ;
      RECT 0 -0.4 1.215 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.15 4.64 15.18 5.44 ;
      RECT 13.81 4.465 14.15 5.44 ;
      RECT 12.53 4.64 13.81 5.44 ;
      RECT 12.19 4.085 12.53 5.44 ;
      RECT 10.465 4.64 12.19 5.44 ;
      RECT 10.125 4.08 10.465 5.44 ;
      RECT 8.37 4.64 10.125 5.44 ;
      RECT 7.43 4.08 8.37 5.44 ;
      RECT 4.07 4.64 7.43 5.44 ;
      RECT 3.73 4.465 4.07 5.44 ;
      RECT 1.48 4.64 3.73 5.44 ;
      RECT 1.14 4.465 1.48 5.44 ;
      RECT 0 4.64 1.14 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.495 1.545 13.725 3.105 ;
      RECT 13.355 1.545 13.495 1.775 ;
      RECT 13.085 2.875 13.495 3.105 ;
      RECT 13.125 1.42 13.355 1.775 ;
      RECT 12.44 2.11 13.1 2.45 ;
      RECT 12.855 2.875 13.085 3.35 ;
      RECT 12.21 1.865 12.44 3.76 ;
      RECT 11.65 1.865 12.21 2.095 ;
      RECT 11.17 3.53 12.21 3.76 ;
      RECT 11.285 0.915 11.65 2.095 ;
      RECT 10.24 3.06 11.535 3.29 ;
      RECT 10.93 1.865 11.285 2.095 ;
      RECT 10.83 3.53 11.17 3.96 ;
      RECT 10.83 1.865 10.93 2.57 ;
      RECT 10.7 1.865 10.83 2.58 ;
      RECT 10.49 2.24 10.7 2.58 ;
      RECT 10.01 1.55 10.24 3.29 ;
      RECT 9.315 1.55 10.01 1.78 ;
      RECT 9.765 3.06 10.01 3.29 ;
      RECT 9.465 3.06 9.765 4.34 ;
      RECT 9.24 2.39 9.47 2.79 ;
      RECT 9.425 4 9.465 4.34 ;
      RECT 9.085 1.29 9.315 1.78 ;
      RECT 8.875 2.56 9.24 2.79 ;
      RECT 8.645 2.56 8.875 3.85 ;
      RECT 8.415 2.09 8.855 2.32 ;
      RECT 7.185 3.62 8.645 3.85 ;
      RECT 8.185 0.675 8.415 3.385 ;
      RECT 6.745 0.675 8.185 0.905 ;
      RECT 7.43 3.155 8.185 3.385 ;
      RECT 7.685 2.305 7.915 2.67 ;
      RECT 6.725 2.305 7.685 2.56 ;
      RECT 6.955 2.81 7.185 4.365 ;
      RECT 4.53 4.135 6.955 4.365 ;
      RECT 6.405 0.635 6.745 0.975 ;
      RECT 6.495 1.825 6.725 3.69 ;
      RECT 5.705 1.825 6.495 2.055 ;
      RECT 5.75 3.46 6.495 3.69 ;
      RECT 5.925 2.44 6.265 2.78 ;
      RECT 5.015 2.495 5.925 2.725 ;
      RECT 5.41 3.46 5.75 3.8 ;
      RECT 5.475 1.1 5.705 2.055 ;
      RECT 3.875 1.655 5.475 1.885 ;
      RECT 5.12 0.77 5.23 1.11 ;
      RECT 4.89 0.77 5.12 1.42 ;
      RECT 4.99 2.115 5.015 2.725 ;
      RECT 4.76 2.115 4.99 3.87 ;
      RECT 3.305 1.19 4.89 1.42 ;
      RECT 4.675 2.115 4.76 2.455 ;
      RECT 4.3 4.005 4.53 4.365 ;
      RECT 3.345 4.005 4.3 4.235 ;
      RECT 3.535 1.655 3.875 2.08 ;
      RECT 3.115 4.005 3.345 4.32 ;
      RECT 3.075 1.19 3.305 3.605 ;
      RECT 2.325 4.09 3.115 4.32 ;
      RECT 2.915 1.19 3.075 1.42 ;
      RECT 2.785 3.375 3.075 3.605 ;
      RECT 2.575 0.965 2.915 1.42 ;
      RECT 2.555 3.375 2.785 3.8 ;
      RECT 2.35 1.89 2.58 3.06 ;
      RECT 2.325 2.83 2.35 3.06 ;
      RECT 2.095 2.83 2.325 4.32 ;
      RECT 2.075 3.995 2.095 4.32 ;
      RECT 0.765 3.995 2.075 4.225 ;
      RECT 0.6 1.11 0.94 1.45 ;
      RECT 0.545 3.515 0.765 4.225 ;
      RECT 0.545 1.22 0.6 1.45 ;
      RECT 0.315 1.22 0.545 4.225 ;
  END
END DFFRXL

MACRO DFFRX4
  CLASS CORE ;
  FOREIGN DFFRX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 19.8 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4068 ;
  ANTENNAPARTIALMETALAREA 0.345 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.02 2.745 4.48 3.495 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2718 ;
  ANTENNAPARTIALMETALAREA 0.7831 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5917 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.3 1.195 17.68 3.22 ;
      RECT 17.28 1.195 17.3 1.535 ;
      RECT 17.28 2.78 17.3 3.12 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2718 ;
  ANTENNAPARTIALMETALAREA 0.7685 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5705 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.9 1.26 19 3.12 ;
      RECT 18.62 1.195 18.9 3.12 ;
      RECT 18.615 1.195 18.62 2.075 ;
      RECT 18.56 2.78 18.62 3.12 ;
      RECT 18.56 1.195 18.615 1.535 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.198 ;
  ANTENNAPARTIALMETALAREA 0.2457 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0653 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.425 2.71 1.845 3.295 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2844 ;
  ANTENNAPARTIALMETALAREA 0.3523 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3197 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.745 1.85 1.18 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.54 -0.4 19.8 0.4 ;
      RECT 19.2 -0.4 19.54 0.95 ;
      RECT 18.26 -0.4 19.2 0.4 ;
      RECT 17.92 -0.4 18.26 0.95 ;
      RECT 16.98 -0.4 17.92 0.4 ;
      RECT 16.64 -0.4 16.98 0.95 ;
      RECT 15.61 -0.4 16.64 0.4 ;
      RECT 15.27 -0.4 15.61 0.95 ;
      RECT 14.17 -0.4 15.27 0.4 ;
      RECT 13.83 -0.4 14.17 0.95 ;
      RECT 12.71 -0.4 13.83 0.4 ;
      RECT 12.37 -0.4 12.71 0.95 ;
      RECT 10.94 -0.4 12.37 0.4 ;
      RECT 10.6 -0.4 10.94 1.08 ;
      RECT 8.345 -0.4 10.6 0.4 ;
      RECT 8.115 -0.4 8.345 1.475 ;
      RECT 6.49 -0.4 8.115 0.4 ;
      RECT 7.93 1.245 8.115 1.475 ;
      RECT 6.15 -0.4 6.49 0.96 ;
      RECT 4.865 -0.4 6.15 0.4 ;
      RECT 4.525 -0.4 4.865 1.335 ;
      RECT 1.295 -0.4 4.525 0.4 ;
      RECT 0.955 -0.4 1.295 0.575 ;
      RECT 0 -0.4 0.955 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.54 4.64 19.8 5.44 ;
      RECT 19.2 4.04 19.54 5.44 ;
      RECT 18.26 4.64 19.2 5.44 ;
      RECT 17.92 4.04 18.26 5.44 ;
      RECT 16.98 4.64 17.92 5.44 ;
      RECT 16.64 4.04 16.98 5.44 ;
      RECT 15.41 4.64 16.64 5.44 ;
      RECT 15.07 2.845 15.41 5.44 ;
      RECT 12.81 4.64 15.07 5.44 ;
      RECT 12.47 4.08 12.81 5.44 ;
      RECT 10.33 4.64 12.47 5.44 ;
      RECT 9.99 3.675 10.33 5.44 ;
      RECT 7.48 4.64 9.99 5.44 ;
      RECT 7.14 3.92 7.48 5.44 ;
      RECT 3.82 4.64 7.14 5.44 ;
      RECT 3.48 4.465 3.82 5.44 ;
      RECT 1.545 4.64 3.48 5.44 ;
      RECT 1.15 4.385 1.545 5.44 ;
      RECT 0 4.64 1.15 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 19.305 2.03 19.535 3.75 ;
      RECT 16.975 3.52 19.305 3.75 ;
      RECT 16.745 1.395 16.975 3.75 ;
      RECT 16.29 1.395 16.745 1.73 ;
      RECT 16.13 3.265 16.745 3.495 ;
      RECT 15.51 2.1 16.45 2.44 ;
      RECT 15.95 1.39 16.29 1.73 ;
      RECT 15.79 2.975 16.13 3.785 ;
      RECT 15.94 1.395 15.95 1.675 ;
      RECT 14.89 2.155 15.51 2.385 ;
      RECT 14.66 0.72 14.89 2.69 ;
      RECT 14.55 0.72 14.66 1.475 ;
      RECT 14.13 2.46 14.66 2.69 ;
      RECT 13.45 1.245 14.55 1.475 ;
      RECT 14.055 1.725 14.41 2.065 ;
      RECT 13.9 2.46 14.13 3.835 ;
      RECT 13.47 1.725 14.055 2.105 ;
      RECT 13.79 2.985 13.9 3.835 ;
      RECT 12.2 3.605 13.79 3.835 ;
      RECT 12.465 1.875 13.47 2.105 ;
      RECT 13.22 0.7 13.45 1.475 ;
      RECT 13.11 0.7 13.22 1.04 ;
      RECT 12.235 1.495 12.465 3.365 ;
      RECT 9.895 1.495 12.235 1.735 ;
      RECT 11.605 3.135 12.235 3.365 ;
      RECT 11.97 3.605 12.2 4.25 ;
      RECT 11.465 2.425 11.805 2.82 ;
      RECT 11.605 3.75 11.66 4.09 ;
      RECT 11.375 3.135 11.605 4.09 ;
      RECT 9.435 2.425 11.465 2.655 ;
      RECT 9.695 3.135 11.375 3.365 ;
      RECT 11.32 3.75 11.375 4.09 ;
      RECT 9.665 1.105 9.895 1.735 ;
      RECT 9.465 3.135 9.695 3.855 ;
      RECT 9.25 1.105 9.665 1.335 ;
      RECT 9.05 3.625 9.465 3.855 ;
      RECT 9.205 1.75 9.435 2.655 ;
      RECT 8.92 2.425 9.205 2.655 ;
      RECT 8.71 3.625 9.05 3.99 ;
      RECT 8.69 1.745 8.92 3.145 ;
      RECT 7.465 1.745 8.69 1.975 ;
      RECT 8.245 2.915 8.69 3.145 ;
      RECT 6.875 2.235 8.46 2.465 ;
      RECT 8.24 2.915 8.245 3.945 ;
      RECT 8.015 2.915 8.24 4 ;
      RECT 7.9 3.66 8.015 4 ;
      RECT 7.505 2.84 7.67 3.18 ;
      RECT 7.275 2.84 7.505 3.66 ;
      RECT 7.235 0.675 7.465 1.975 ;
      RECT 6.745 3.43 7.275 3.66 ;
      RECT 6.74 0.675 7.235 0.905 ;
      RECT 6.645 1.565 6.875 3.145 ;
      RECT 6.515 3.43 6.745 4.365 ;
      RECT 5.93 1.565 6.645 1.795 ;
      RECT 6.2 2.915 6.645 3.145 ;
      RECT 4.365 4.135 6.515 4.365 ;
      RECT 5.86 2.915 6.2 3.87 ;
      RECT 5.83 2.1 6.17 2.44 ;
      RECT 5.59 1.43 5.93 1.795 ;
      RECT 5.015 2.155 5.83 2.385 ;
      RECT 3.55 1.565 5.59 1.795 ;
      RECT 5.015 3.56 5.07 3.9 ;
      RECT 4.785 2.025 5.015 3.9 ;
      RECT 4.27 2.025 4.785 2.255 ;
      RECT 4.73 3.56 4.785 3.9 ;
      RECT 4.135 3.945 4.365 4.365 ;
      RECT 2.575 0.825 4.275 1.055 ;
      RECT 3.165 3.945 4.135 4.175 ;
      RECT 3.55 2.32 3.66 2.66 ;
      RECT 3.32 1.565 3.55 2.66 ;
      RECT 2.955 3.035 3.165 4.4 ;
      RECT 2.935 1.775 2.955 4.4 ;
      RECT 2.725 1.775 2.935 3.265 ;
      RECT 2.02 4.17 2.935 4.4 ;
      RECT 2.09 1.775 2.725 2.005 ;
      RECT 2.49 3.5 2.62 3.84 ;
      RECT 2.345 0.825 2.575 1.47 ;
      RECT 2.26 2.24 2.49 3.84 ;
      RECT 2.235 1.13 2.345 1.47 ;
      RECT 1.85 2.24 2.26 2.47 ;
      RECT 1.85 1.185 2.235 1.415 ;
      RECT 1.79 3.71 2.02 4.4 ;
      RECT 1.62 1.185 1.85 2.47 ;
      RECT 0.605 3.71 1.79 3.94 ;
      RECT 0.495 1.22 0.635 1.56 ;
      RECT 0.495 3.01 0.605 3.94 ;
      RECT 0.295 1.22 0.495 3.94 ;
      RECT 0.265 1.275 0.295 3.94 ;
  END
END DFFRX4

MACRO DFFRX2
  CLASS CORE ;
  FOREIGN DFFRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.3098 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.605 2.875 4.66 3.39 ;
      RECT 4.32 2.755 4.605 3.39 ;
      RECT 4.175 2.755 4.32 3.335 ;
      RECT 4.13 2.875 4.175 3.24 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1919 ;
  ANTENNAPARTIALMETALAREA 0.7511 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8408 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.57 1.515 15.71 2.13 ;
      RECT 15.565 2.93 15.62 3.27 ;
      RECT 15.565 1.26 15.57 2.13 ;
      RECT 15.335 1.26 15.565 3.27 ;
      RECT 15.15 1.26 15.335 2.13 ;
      RECT 15.28 2.93 15.335 3.27 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1995 ;
  ANTENNAPARTIALMETALAREA 0.6729 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6659 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17 1.26 17.005 3.23 ;
      RECT 16.705 1.26 17 3.275 ;
      RECT 16.64 1.26 16.705 1.6 ;
      RECT 16.57 2.93 16.705 3.275 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3192 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2932 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.935 1.84 3.775 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.3219 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.785 1.26 1.18 2.075 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.28 -0.4 17.16 0.4 ;
      RECT 15.94 -0.4 16.28 0.95 ;
      RECT 14.12 -0.4 15.94 0.4 ;
      RECT 13.78 -0.4 14.12 1.36 ;
      RECT 12.63 -0.4 13.78 0.4 ;
      RECT 12.29 -0.4 12.63 0.575 ;
      RECT 10.77 -0.4 12.29 0.4 ;
      RECT 10.43 -0.4 10.77 1.25 ;
      RECT 8.04 -0.4 10.43 0.4 ;
      RECT 7.7 -0.4 8.04 1.37 ;
      RECT 6.34 -0.4 7.7 0.4 ;
      RECT 6 -0.4 6.34 0.96 ;
      RECT 5.12 -0.4 6 0.44 ;
      RECT 4.695 -0.4 5.12 1.335 ;
      RECT 1.3 -0.4 4.695 0.4 ;
      RECT 0.96 -0.4 1.3 0.575 ;
      RECT 0 -0.4 0.96 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.26 4.64 17.16 5.44 ;
      RECT 15.92 4.08 16.26 5.44 ;
      RECT 14.2 4.64 15.92 5.44 ;
      RECT 13.86 3.68 14.2 5.44 ;
      RECT 11.42 4.64 13.86 5.44 ;
      RECT 11.08 4.08 11.42 5.44 ;
      RECT 8.705 4.64 11.08 5.44 ;
      RECT 7.26 4.135 8.705 5.44 ;
      RECT 4.36 4.64 7.26 5.44 ;
      RECT 4.02 4.465 4.36 5.44 ;
      RECT 1.46 4.64 4.02 5.44 ;
      RECT 1.12 4.465 1.46 5.44 ;
      RECT 0 4.64 1.12 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 16.245 1.91 16.475 2.655 ;
      RECT 16.2 2.425 16.245 2.655 ;
      RECT 15.97 2.425 16.2 3.805 ;
      RECT 14.92 3.575 15.97 3.805 ;
      RECT 14.81 3.575 14.92 4.02 ;
      RECT 14.81 1.02 14.84 1.36 ;
      RECT 14.58 1.02 14.81 4.02 ;
      RECT 14.5 1.02 14.58 1.36 ;
      RECT 14.295 1.63 14.35 2.045 ;
      RECT 14.065 1.63 14.295 3.165 ;
      RECT 14.01 1.63 14.065 2.045 ;
      RECT 13.52 2.935 14.065 3.165 ;
      RECT 13.4 1.815 14.01 2.045 ;
      RECT 13.29 2.935 13.52 3.51 ;
      RECT 13.17 0.91 13.4 2.045 ;
      RECT 12.74 3.28 13.29 3.51 ;
      RECT 13.06 0.91 13.17 1.25 ;
      RECT 12.49 1.815 13.17 2.045 ;
      RECT 12.63 3.28 12.74 3.62 ;
      RECT 12.4 3.28 12.63 4.27 ;
      RECT 12.05 2.46 12.55 2.8 ;
      RECT 12.205 1.63 12.49 2.045 ;
      RECT 12.12 3.93 12.4 4.27 ;
      RECT 12.15 1.63 12.205 1.97 ;
      RECT 11.92 2.46 12.05 3.335 ;
      RECT 11.69 1.685 11.92 3.335 ;
      RECT 11.59 1.685 11.69 1.915 ;
      RECT 11.68 2.68 11.69 3.335 ;
      RECT 10.665 3.105 11.68 3.335 ;
      RECT 11.36 1.225 11.59 1.915 ;
      RECT 11.405 2.205 11.46 2.435 ;
      RECT 11.175 2.205 11.405 2.44 ;
      RECT 11.13 1.225 11.36 1.755 ;
      RECT 10.785 2.21 11.175 2.44 ;
      RECT 9.46 1.525 11.13 1.755 ;
      RECT 10.555 1.985 10.785 2.44 ;
      RECT 10.435 3.105 10.665 3.48 ;
      RECT 9 1.985 10.555 2.215 ;
      RECT 10.1 3.25 10.435 3.48 ;
      RECT 9.76 3.25 10.1 3.59 ;
      RECT 9.52 2.6 9.86 2.94 ;
      RECT 9.505 2.71 9.52 2.94 ;
      RECT 9.275 2.71 9.505 3.9 ;
      RECT 9.23 1.09 9.46 1.755 ;
      RECT 7.375 3.67 9.275 3.9 ;
      RECT 9.06 1.09 9.23 1.43 ;
      RECT 8.77 1.705 9 3.44 ;
      RECT 7.24 1.705 8.77 1.935 ;
      RECT 7.83 3.21 8.77 3.44 ;
      RECT 8.2 2.17 8.54 2.885 ;
      RECT 6.575 2.17 8.2 2.4 ;
      RECT 7.53 2.63 7.87 2.97 ;
      RECT 7.375 2.685 7.53 2.97 ;
      RECT 7.145 2.685 7.375 3.9 ;
      RECT 7.235 1.205 7.24 1.935 ;
      RECT 7.125 1.15 7.235 1.935 ;
      RECT 6.935 3.67 7.145 3.9 ;
      RECT 6.95 0.665 7.125 1.935 ;
      RECT 6.895 0.665 6.95 1.49 ;
      RECT 6.705 3.67 6.935 4.355 ;
      RECT 6.63 0.665 6.895 0.895 ;
      RECT 4.825 4.125 6.705 4.355 ;
      RECT 6.345 1.575 6.575 3.185 ;
      RECT 5.84 1.575 6.345 1.805 ;
      RECT 6.155 2.955 6.345 3.185 ;
      RECT 6.155 3.47 6.21 3.81 ;
      RECT 5.925 2.955 6.155 3.81 ;
      RECT 5.775 2.14 6.115 2.48 ;
      RECT 5.87 3.47 5.925 3.81 ;
      RECT 5.61 1.455 5.84 1.805 ;
      RECT 5.345 2.195 5.775 2.425 ;
      RECT 5.5 1.455 5.61 1.795 ;
      RECT 3.68 1.565 5.5 1.795 ;
      RECT 5.345 3.55 5.4 3.89 ;
      RECT 5.115 2.195 5.345 3.89 ;
      RECT 5.11 2.195 5.115 2.425 ;
      RECT 5.06 3.55 5.115 3.89 ;
      RECT 4.56 2.03 5.11 2.425 ;
      RECT 4.595 3.945 4.825 4.355 ;
      RECT 3.705 3.945 4.595 4.175 ;
      RECT 4.08 0.675 4.42 1.11 ;
      RECT 3.025 0.675 4.08 0.905 ;
      RECT 3.475 3.945 3.705 4.255 ;
      RECT 3.35 1.565 3.68 2.085 ;
      RECT 2.56 4.025 3.475 4.255 ;
      RECT 3.34 1.745 3.35 2.085 ;
      RECT 3.045 3.3 3.1 3.64 ;
      RECT 3.025 3.28 3.045 3.64 ;
      RECT 2.795 0.675 3.025 3.64 ;
      RECT 2.43 0.675 2.795 1.27 ;
      RECT 2.76 3.3 2.795 3.64 ;
      RECT 2.46 3.97 2.56 4.31 ;
      RECT 2.415 1.59 2.46 4.31 ;
      RECT 2.375 0.905 2.43 1.27 ;
      RECT 2.23 1.535 2.415 4.31 ;
      RECT 2.32 0.93 2.375 1.27 ;
      RECT 2.075 1.535 2.23 1.875 ;
      RECT 2.22 3.97 2.23 4.31 ;
      RECT 0.5 4.005 2.22 4.235 ;
      RECT 0.5 1.105 0.555 1.445 ;
      RECT 0.5 3.055 0.555 3.395 ;
      RECT 0.27 1.105 0.5 4.235 ;
      RECT 0.215 1.105 0.27 1.445 ;
      RECT 0.215 3.055 0.27 3.395 ;
  END
END DFFRX2

MACRO DFFRX1
  CLASS CORE ;
  FOREIGN DFFRX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.18 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.332 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4257 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.525 3.34 4.825 3.57 ;
      RECT 4.13 2.95 4.525 3.57 ;
      RECT 4.1 2.965 4.13 3.57 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6496 ;
  ANTENNAPARTIALMETALAREA 1.0749 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9555 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.18 2.035 14.41 3.295 ;
      RECT 13.575 2.035 14.18 2.265 ;
      RECT 13.89 3.065 14.18 3.295 ;
      RECT 13.66 3.065 13.89 3.795 ;
      RECT 13.52 3.5 13.66 3.795 ;
      RECT 13.345 1.38 13.575 2.265 ;
      RECT 13.18 3.5 13.52 3.99 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.8519 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5722 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.78 1.27 14.995 3.93 ;
      RECT 14.735 1.27 14.78 3.98 ;
      RECT 14.66 1.27 14.735 1.845 ;
      RECT 14.44 3.64 14.735 3.98 ;
      RECT 14.63 1.355 14.66 1.845 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2825 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.635 2.94 1.84 3.305 ;
      RECT 1.3 2.69 1.635 3.305 ;
      RECT 1.295 2.69 1.3 3.03 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.2541 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 1.775 1.185 2.435 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.29 -0.4 15.18 0.4 ;
      RECT 13.95 -0.4 14.29 0.575 ;
      RECT 12.21 -0.4 13.95 0.4 ;
      RECT 11.87 -0.4 12.21 0.575 ;
      RECT 10.69 -0.4 11.87 0.4 ;
      RECT 10.35 -0.4 10.69 1.31 ;
      RECT 6.035 -0.4 10.35 0.4 ;
      RECT 7.81 1.44 7.92 1.78 ;
      RECT 7.58 1.205 7.81 1.78 ;
      RECT 6.33 1.205 7.58 1.435 ;
      RECT 6.035 1.205 6.33 1.525 ;
      RECT 5.805 -0.4 6.035 1.525 ;
      RECT 4.19 -0.4 5.805 0.4 ;
      RECT 3.85 -0.4 4.19 0.96 ;
      RECT 1.46 -0.4 3.85 0.4 ;
      RECT 1.12 -0.4 1.46 0.575 ;
      RECT 0 -0.4 1.12 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.1 4.64 15.18 5.44 ;
      RECT 13.76 4.465 14.1 5.44 ;
      RECT 12.76 4.64 13.76 5.44 ;
      RECT 12.42 3.62 12.76 5.44 ;
      RECT 10.74 4.64 12.42 5.44 ;
      RECT 10.4 4.07 10.74 5.44 ;
      RECT 8.4 4.64 10.4 5.44 ;
      RECT 7.46 4.07 8.4 5.44 ;
      RECT 4.33 4.64 7.46 5.44 ;
      RECT 3.99 4.465 4.33 5.44 ;
      RECT 1.605 4.64 3.99 5.44 ;
      RECT 1.195 4.39 1.605 5.44 ;
      RECT 0 4.64 1.195 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.42 2.495 13.95 2.835 ;
      RECT 13.1 2.495 13.42 3.14 ;
      RECT 13.08 1.25 13.1 3.14 ;
      RECT 12.8 1.25 13.08 2.795 ;
      RECT 12.77 1.25 12.8 1.55 ;
      RECT 12.43 1.21 12.77 1.55 ;
      RECT 12.455 1.825 12.56 2.11 ;
      RECT 12.225 1.825 12.455 3.295 ;
      RECT 11.925 1.825 12.225 2.055 ;
      RECT 11.48 3.065 12.225 3.295 ;
      RECT 11.695 1.595 11.925 2.055 ;
      RECT 11.39 1.595 11.695 1.825 ;
      RECT 11.14 3.065 11.48 3.94 ;
      RECT 11.39 0.97 11.45 1.31 ;
      RECT 11.11 0.97 11.39 1.825 ;
      RECT 11.325 2.14 11.38 2.48 ;
      RECT 11.04 2.14 11.325 2.505 ;
      RECT 10.54 1.595 11.11 1.825 ;
      RECT 9.915 2.275 11.04 2.505 ;
      RECT 10.255 1.595 10.54 2.045 ;
      RECT 10.2 1.705 10.255 2.045 ;
      RECT 9.915 4 10.03 4.34 ;
      RECT 9.905 2.275 9.915 4.34 ;
      RECT 9.685 1.285 9.905 4.34 ;
      RECT 9.675 1.285 9.685 4.285 ;
      RECT 9.28 1.285 9.675 1.515 ;
      RECT 8.94 1.23 9.28 1.57 ;
      RECT 9.15 2.5 9.26 2.84 ;
      RECT 8.92 2.5 9.15 3.84 ;
      RECT 7.525 3.61 8.92 3.84 ;
      RECT 8.535 1.83 8.915 2.17 ;
      RECT 8.305 0.675 8.535 3.375 ;
      RECT 6.605 0.675 8.305 0.905 ;
      RECT 7.76 3.145 8.305 3.375 ;
      RECT 8.005 2.02 8.06 2.41 ;
      RECT 7.72 2.02 8.005 2.415 ;
      RECT 6.645 2.18 7.72 2.415 ;
      RECT 7.295 2.705 7.525 3.84 ;
      RECT 7.165 3.61 7.295 3.84 ;
      RECT 6.935 3.61 7.165 4.365 ;
      RECT 4.79 4.135 6.935 4.365 ;
      RECT 6.415 1.825 6.645 3.385 ;
      RECT 6.265 0.635 6.605 0.975 ;
      RECT 5.575 1.825 6.415 2.055 ;
      RECT 6.11 3.155 6.415 3.385 ;
      RECT 5.88 3.155 6.11 3.82 ;
      RECT 5.76 2.44 6.1 2.78 ;
      RECT 5.77 3.48 5.88 3.82 ;
      RECT 5.355 2.495 5.76 2.725 ;
      RECT 5.37 1.655 5.575 2.055 ;
      RECT 5.355 3.48 5.41 3.82 ;
      RECT 5.345 1.14 5.37 2.055 ;
      RECT 5.125 2.435 5.355 3.82 ;
      RECT 5.14 1.14 5.345 1.885 ;
      RECT 3.825 1.655 5.14 1.885 ;
      RECT 4.99 2.435 5.125 2.665 ;
      RECT 5.07 3.48 5.125 3.82 ;
      RECT 4.6 2.115 4.99 2.665 ;
      RECT 4.755 0.77 4.87 1.11 ;
      RECT 4.56 3.945 4.79 4.365 ;
      RECT 4.525 0.77 4.755 1.42 ;
      RECT 3.675 3.945 4.56 4.175 ;
      RECT 2.825 1.19 4.525 1.42 ;
      RECT 3.485 1.655 3.825 2.08 ;
      RECT 3.465 2.935 3.675 4.355 ;
      RECT 3.445 2.395 3.465 4.355 ;
      RECT 3.235 2.395 3.445 3.165 ;
      RECT 2.155 4.125 3.445 4.355 ;
      RECT 2.905 2.395 3.235 2.625 ;
      RECT 2.775 3.48 3.11 3.84 ;
      RECT 2.675 1.995 2.905 2.625 ;
      RECT 2.485 1.16 2.825 1.5 ;
      RECT 2.545 2.965 2.775 3.84 ;
      RECT 2.335 1.995 2.675 2.225 ;
      RECT 2.37 2.965 2.545 3.195 ;
      RECT 2.1 1.27 2.485 1.5 ;
      RECT 2.14 2.46 2.37 3.195 ;
      RECT 1.925 3.745 2.155 4.355 ;
      RECT 2.1 2.46 2.14 2.69 ;
      RECT 1.87 1.27 2.1 2.69 ;
      RECT 0.6 3.745 1.925 3.975 ;
      RECT 0.545 1.1 0.85 1.44 ;
      RECT 0.545 3.52 0.6 3.975 ;
      RECT 0.315 1.1 0.545 3.975 ;
      RECT 0.26 3.52 0.315 3.975 ;
  END
END DFFRX1

MACRO DFFNSRXL
  CLASS CORE ;
  FOREIGN DFFNSRXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.288 ;
  ANTENNAPARTIALMETALAREA 1.7841 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.427 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.555 4.075 11.665 4.365 ;
      RECT 11.325 4.02 11.555 4.365 ;
      RECT 8.795 4.135 11.325 4.365 ;
      RECT 8.37 4.125 8.795 4.365 ;
      RECT 5.875 4.125 8.37 4.355 ;
      RECT 5.645 4.005 5.875 4.355 ;
      RECT 4.695 4.005 5.645 4.235 ;
      RECT 4.465 4.005 4.695 4.365 ;
      RECT 4.32 4.135 4.465 4.365 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2225 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.98 1.765 6.4 2.295 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5792 ;
  ANTENNAPARTIALMETALAREA 0.6996 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1535 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.215 1.095 15.37 1.435 ;
      RECT 14.985 1.095 15.215 3.4 ;
      RECT 14.735 2.965 14.985 3.4 ;
      RECT 14.7 3.17 14.735 3.4 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.576 ;
  ANTENNAPARTIALMETALAREA 0.7264 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3231 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.835 2.955 16.945 3.195 ;
      RECT 16.77 1.095 16.835 3.195 ;
      RECT 16.605 1.095 16.77 3.58 ;
      RECT 16.47 1.095 16.605 1.435 ;
      RECT 16.43 2.965 16.605 3.58 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.4083 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5635 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 1.72 1.18 2.62 ;
      RECT 0.605 2.28 0.8 2.62 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0017 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.14 1.885 2.66 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.09 -0.4 17.16 0.4 ;
      RECT 15.75 -0.4 16.09 1.435 ;
      RECT 14.53 -0.4 15.75 0.4 ;
      RECT 14.19 -0.4 14.53 0.575 ;
      RECT 11.335 -0.4 14.19 0.4 ;
      RECT 10.995 -0.4 11.335 0.575 ;
      RECT 8.77 -0.4 10.995 0.4 ;
      RECT 8.43 -0.4 8.77 1.43 ;
      RECT 7.005 -0.4 8.43 0.4 ;
      RECT 6.775 -0.4 7.005 0.9 ;
      RECT 4.105 -0.4 6.775 0.4 ;
      RECT 3.765 -0.4 4.105 0.9 ;
      RECT 1.425 -0.4 3.765 0.4 ;
      RECT 1.085 -0.4 1.425 0.575 ;
      RECT 0 -0.4 1.085 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.95 4.64 17.16 5.44 ;
      RECT 15.61 4.09 15.95 5.44 ;
      RECT 13.45 4.64 15.61 5.44 ;
      RECT 13.11 3.395 13.45 5.44 ;
      RECT 12.285 4.64 13.11 5.44 ;
      RECT 12.055 3.395 12.285 5.44 ;
      RECT 11.37 3.395 12.055 3.625 ;
      RECT 5.415 4.64 12.055 5.44 ;
      RECT 11.01 3.31 11.37 3.625 ;
      RECT 10.785 3.395 11.01 3.625 ;
      RECT 10.555 3.395 10.785 3.845 ;
      RECT 8.845 3.615 10.555 3.845 ;
      RECT 8.615 3.515 8.845 3.845 ;
      RECT 8.375 3.515 8.615 3.745 ;
      RECT 5.075 4.465 5.415 5.44 ;
      RECT 4.09 4.64 5.075 5.44 ;
      RECT 3.75 4.465 4.09 5.44 ;
      RECT 1.1 4.64 3.75 5.44 ;
      RECT 0.76 4.465 1.1 5.44 ;
      RECT 0 4.64 0.76 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.86 2.145 16.33 2.375 ;
      RECT 15.63 2.145 15.86 3.86 ;
      RECT 14.43 3.63 15.63 3.86 ;
      RECT 14.43 1.17 14.54 1.51 ;
      RECT 14.2 1.17 14.43 3.86 ;
      RECT 13.83 3.395 14.2 3.735 ;
      RECT 13.645 1.825 13.875 3.165 ;
      RECT 13.485 0.98 13.735 1.32 ;
      RECT 13.025 1.825 13.645 2.055 ;
      RECT 11.89 2.935 13.645 3.165 ;
      RECT 13.395 0.63 13.485 1.32 ;
      RECT 13.255 0.63 13.395 1.265 ;
      RECT 12.155 0.63 13.255 0.86 ;
      RECT 12.795 1.09 13.025 2.055 ;
      RECT 12.595 1.09 12.795 1.32 ;
      RECT 12.07 1.855 12.3 2.23 ;
      RECT 12.135 0.63 12.155 1.235 ;
      RECT 11.925 0.63 12.135 1.29 ;
      RECT 10.945 1.855 12.07 2.085 ;
      RECT 11.795 0.95 11.925 1.29 ;
      RECT 11.66 2.615 11.89 3.165 ;
      RECT 10.835 2.615 11.66 2.845 ;
      RECT 10.715 1.25 10.945 2.085 ;
      RECT 10.295 1.25 10.715 1.48 ;
      RECT 9.425 0.72 10.585 0.95 ;
      RECT 10.065 1.25 10.295 3.36 ;
      RECT 9.995 1.25 10.065 1.535 ;
      RECT 9.655 3.13 10.065 3.36 ;
      RECT 9.765 1.195 9.995 1.535 ;
      RECT 9.425 2.485 9.75 2.715 ;
      RECT 9.195 0.72 9.425 3.28 ;
      RECT 7.915 1.66 9.195 1.89 ;
      RECT 7.94 3.05 9.195 3.28 ;
      RECT 8.635 2.125 8.865 2.605 ;
      RECT 7.455 2.125 8.635 2.355 ;
      RECT 7.47 2.59 8.225 2.82 ;
      RECT 7.71 3.05 7.94 3.8 ;
      RECT 7.685 0.67 7.915 1.89 ;
      RECT 7.475 0.67 7.685 0.9 ;
      RECT 7.24 2.59 7.47 3.84 ;
      RECT 7.225 1.135 7.455 2.355 ;
      RECT 6.335 3.61 7.24 3.84 ;
      RECT 5.745 1.135 7.225 1.365 ;
      RECT 6.755 1.635 6.985 3.375 ;
      RECT 6.57 2.805 6.755 3.375 ;
      RECT 5.595 2.805 6.57 3.035 ;
      RECT 6.105 3.535 6.335 3.84 ;
      RECT 3.325 3.535 6.105 3.765 ;
      RECT 5.515 1.135 5.745 2.575 ;
      RECT 5.505 1.135 5.515 1.435 ;
      RECT 5.31 2.345 5.515 2.575 ;
      RECT 5.165 1.095 5.505 1.435 ;
      RECT 5.08 2.345 5.31 3.305 ;
      RECT 4.55 1.695 5.225 1.925 ;
      RECT 4.065 3.075 5.08 3.305 ;
      RECT 4.32 1.6 4.55 1.925 ;
      RECT 3.6 1.6 4.32 1.83 ;
      RECT 3.835 2.065 4.065 3.305 ;
      RECT 3.595 1.3 3.6 1.83 ;
      RECT 3.365 1.29 3.595 2.965 ;
      RECT 2.935 1.29 3.365 1.53 ;
      RECT 2.835 2.735 3.365 2.965 ;
      RECT 3.095 3.535 3.325 4.28 ;
      RECT 2.35 1.77 3.12 2.11 ;
      RECT 2.355 4.05 3.095 4.28 ;
      RECT 2.65 0.9 2.935 1.53 ;
      RECT 2.605 2.735 2.835 3.82 ;
      RECT 2.595 0.9 2.65 1.24 ;
      RECT 2.35 2.93 2.355 4.28 ;
      RECT 2.125 1.505 2.35 4.28 ;
      RECT 1.785 0.675 2.17 1.04 ;
      RECT 2.12 1.505 2.125 3.48 ;
      RECT 2.075 1.505 2.12 1.79 ;
      RECT 1.995 3.02 2.12 3.48 ;
      RECT 1.735 1.45 2.075 1.79 ;
      RECT 1.52 3.02 1.995 3.25 ;
      RECT 1.48 3.835 1.805 4.39 ;
      RECT 0.465 0.81 1.785 1.04 ;
      RECT 0.48 3.835 1.48 4.065 ;
      RECT 0.48 2.925 0.535 3.265 ;
      RECT 0.25 2.925 0.48 4.065 ;
      RECT 0.235 0.81 0.465 1.77 ;
      RECT 0.195 2.925 0.25 3.265 ;
  END
END DFFNSRXL

MACRO DFFNSRX4
  CLASS CORE ;
  FOREIGN DFFNSRX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 23.1 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9792 ;
  ANTENNAPARTIALMETALAREA 2.2402 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.5682 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.73 4 14.32 4.23 ;
      RECT 8.5 4 8.73 4.29 ;
      RECT 8.365 4.06 8.5 4.29 ;
      RECT 8.135 4.06 8.365 4.335 ;
      RECT 4.685 4.105 8.135 4.335 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4461 ;
  ANTENNAPARTIALMETALAREA 0.2326 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.595 2.295 7.065 2.79 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2857 ;
  ANTENNAPARTIALMETALAREA 0.6799 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.3532 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.98 1.42 21 1.85 ;
      RECT 20.98 2.63 21 3.195 ;
      RECT 20.66 1.42 20.98 3.22 ;
      RECT 20.6 1.82 20.66 3.22 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2857 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.3108 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.28 1.82 22.3 3.22 ;
      RECT 21.94 1.42 22.28 3.22 ;
      RECT 21.92 1.82 21.94 3.22 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2412 ;
  ANTENNAPARTIALMETALAREA 0.2531 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.175 0.555 2.785 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.306 ;
  ANTENNAPARTIALMETALAREA 0.2836 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 2.035 1.49 2.325 ;
      RECT 0.8 1.815 1.18 2.325 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 22.92 -0.4 23.1 0.4 ;
      RECT 22.58 -0.4 22.92 1.03 ;
      RECT 21.64 -0.4 22.58 0.4 ;
      RECT 21.3 -0.4 21.64 1.045 ;
      RECT 20.36 -0.4 21.3 0.4 ;
      RECT 20.02 -0.4 20.36 1.03 ;
      RECT 15.15 -0.4 20.02 0.4 ;
      RECT 14.81 -0.4 15.15 1.05 ;
      RECT 12.265 -0.4 14.81 0.4 ;
      RECT 11.925 -0.4 12.265 1.175 ;
      RECT 9.57 -0.4 11.925 0.4 ;
      RECT 9.34 -0.4 9.57 0.885 ;
      RECT 7.09 -0.4 9.34 0.4 ;
      RECT 6.72 -0.4 7.09 0.83 ;
      RECT 4.335 -0.4 6.72 0.4 ;
      RECT 3.995 -0.4 4.335 0.845 ;
      RECT 1.105 -0.4 3.995 0.4 ;
      RECT 0.765 -0.4 1.105 0.575 ;
      RECT 0 -0.4 0.765 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 22.92 4.64 23.1 5.44 ;
      RECT 22.58 4.035 22.92 5.44 ;
      RECT 21.64 4.64 22.58 5.44 ;
      RECT 21.3 4.035 21.64 5.44 ;
      RECT 20.36 4.64 21.3 5.44 ;
      RECT 20.02 4.035 20.36 5.44 ;
      RECT 17.61 4.64 20.02 5.44 ;
      RECT 17.27 3.64 17.61 5.44 ;
      RECT 15.55 4.64 17.27 5.44 ;
      RECT 15.32 2.92 15.55 5.44 ;
      RECT 13.345 4.64 15.32 5.44 ;
      RECT 13.005 4.465 13.345 5.44 ;
      RECT 12.19 4.64 13.005 5.44 ;
      RECT 11.85 4.465 12.19 5.44 ;
      RECT 9.525 4.64 11.85 5.44 ;
      RECT 9.185 4.465 9.525 5.44 ;
      RECT 4.41 4.64 9.185 5.44 ;
      RECT 4.07 4.465 4.41 5.44 ;
      RECT 1.085 4.64 4.07 5.44 ;
      RECT 0.745 4.465 1.085 5.44 ;
      RECT 0 4.64 0.745 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 22.605 2.21 22.835 3.74 ;
      RECT 20.295 3.51 22.605 3.74 ;
      RECT 20.065 1.67 20.295 3.74 ;
      RECT 19.545 1.67 20.065 1.9 ;
      RECT 19.26 3.4 20.065 3.74 ;
      RECT 19.065 2.16 19.75 2.5 ;
      RECT 19.315 1.44 19.545 1.9 ;
      RECT 18.9 1.375 19.065 3.015 ;
      RECT 18.835 1.375 18.9 3.61 ;
      RECT 18.05 1.375 18.835 1.605 ;
      RECT 18.67 2.785 18.835 3.61 ;
      RECT 18.485 0.675 18.715 1.03 ;
      RECT 18.56 3.085 18.67 3.61 ;
      RECT 18.37 1.86 18.6 2.26 ;
      RECT 16.33 3.085 18.56 3.315 ;
      RECT 17.33 0.675 18.485 0.905 ;
      RECT 16.11 1.86 18.37 2.09 ;
      RECT 17.68 1.205 18.05 1.605 ;
      RECT 16.705 1.375 17.68 1.605 ;
      RECT 16.99 0.675 17.33 1.05 ;
      RECT 15.875 0.675 16.99 0.905 ;
      RECT 16.475 1.14 16.705 1.605 ;
      RECT 16.265 1.14 16.475 1.37 ;
      RECT 16.22 3.085 16.33 3.6 ;
      RECT 15.99 2.455 16.22 3.6 ;
      RECT 15.825 1.86 16.11 2.155 ;
      RECT 14.83 2.455 15.99 2.685 ;
      RECT 15.765 0.675 15.875 1.29 ;
      RECT 13.68 1.925 15.825 2.155 ;
      RECT 15.645 0.675 15.765 1.605 ;
      RECT 15.535 0.95 15.645 1.605 ;
      RECT 14.375 1.375 15.535 1.605 ;
      RECT 14.755 3.535 14.985 4.41 ;
      RECT 14.6 2.455 14.83 3.305 ;
      RECT 8.195 3.535 14.755 3.765 ;
      RECT 12.755 3.075 14.6 3.305 ;
      RECT 14.145 0.97 14.375 1.605 ;
      RECT 13.45 0.875 13.68 2.155 ;
      RECT 13.285 0.875 13.45 1.105 ;
      RECT 13.29 1.925 13.45 2.155 ;
      RECT 13.06 1.925 13.29 2.845 ;
      RECT 11.52 1.405 13.22 1.635 ;
      RECT 11.055 1.925 13.06 2.155 ;
      RECT 12.525 2.385 12.755 3.305 ;
      RECT 12.32 2.385 12.525 2.615 ;
      RECT 11.29 0.675 11.52 1.635 ;
      RECT 10.28 0.675 11.29 0.905 ;
      RECT 10.89 1.755 11.055 3.135 ;
      RECT 10.825 1.22 10.89 3.135 ;
      RECT 10.66 1.22 10.825 1.985 ;
      RECT 10.515 2.905 10.825 3.135 ;
      RECT 10.28 2.3 10.59 2.53 ;
      RECT 10.05 0.675 10.28 3.195 ;
      RECT 8.66 2.965 10.05 3.195 ;
      RECT 9.53 1.53 9.76 2.325 ;
      RECT 9.11 1.53 9.53 1.76 ;
      RECT 8.88 0.935 9.11 1.76 ;
      RECT 7.735 0.935 8.88 1.165 ;
      RECT 8.56 2.565 8.66 3.195 ;
      RECT 8.56 1.4 8.65 2 ;
      RECT 8.43 1.4 8.56 3.195 ;
      RECT 8.42 1.4 8.43 2.795 ;
      RECT 8.33 1.765 8.42 2.795 ;
      RECT 7.965 3.085 8.195 3.765 ;
      RECT 7.605 3.085 7.965 3.315 ;
      RECT 7.605 1.53 7.78 1.76 ;
      RECT 7.505 0.935 7.735 1.295 ;
      RECT 7.68 3.605 7.735 3.835 ;
      RECT 7.45 3.605 7.68 3.84 ;
      RECT 7.375 1.53 7.605 3.315 ;
      RECT 5.695 1.065 7.505 1.295 ;
      RECT 3.83 3.61 7.45 3.84 ;
      RECT 6.17 3.085 7.375 3.315 ;
      RECT 5.94 2.28 6.17 3.315 ;
      RECT 5.465 1.065 5.695 3.375 ;
      RECT 5.4 1.065 5.465 1.435 ;
      RECT 4.13 3.145 5.465 3.375 ;
      RECT 5.005 1.755 5.235 2.24 ;
      RECT 4.755 1.755 5.005 1.985 ;
      RECT 4.525 1.565 4.755 1.985 ;
      RECT 3.6 1.565 4.525 1.795 ;
      RECT 3.9 2.33 4.13 3.375 ;
      RECT 3.6 3.61 3.83 4.41 ;
      RECT 3.37 0.785 3.6 3.08 ;
      RECT 2.835 4.18 3.6 4.41 ;
      RECT 2.84 0.785 3.37 1.015 ;
      RECT 3.3 2.85 3.37 3.08 ;
      RECT 3.07 2.85 3.3 3.825 ;
      RECT 3.08 1.75 3.135 2.09 ;
      RECT 2.795 1.75 3.08 2.1 ;
      RECT 2.605 2.905 2.835 4.41 ;
      RECT 1.975 1.755 2.795 2.1 ;
      RECT 1.975 2.905 2.605 3.135 ;
      RECT 2.265 0.725 2.46 0.955 ;
      RECT 2.055 3.735 2.37 4.17 ;
      RECT 2.035 0.725 2.265 1.045 ;
      RECT 0.52 3.82 2.055 4.05 ;
      RECT 0.545 0.815 2.035 1.045 ;
      RECT 1.745 1.425 1.975 3.36 ;
      RECT 1.565 1.425 1.745 1.655 ;
      RECT 1.525 3.02 1.745 3.36 ;
      RECT 0.315 0.815 0.545 1.635 ;
      RECT 0.29 3.21 0.52 4.05 ;
      RECT 0.205 1.295 0.315 1.635 ;
      RECT 0.18 3.21 0.29 3.55 ;
  END
END DFFNSRX4

MACRO DFFNSRX2
  CLASS CORE ;
  FOREIGN DFFNSRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5328 ;
  ANTENNAPARTIALMETALAREA 1.8156 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.3422 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.23 3.995 11.74 4.365 ;
      RECT 11.005 4.085 11.23 4.365 ;
      RECT 8.795 4.135 11.005 4.365 ;
      RECT 8.37 4.125 8.795 4.365 ;
      RECT 5.845 4.125 8.37 4.355 ;
      RECT 5.615 4.005 5.845 4.355 ;
      RECT 4.765 4.005 5.615 4.235 ;
      RECT 4.425 4.005 4.765 4.29 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2741 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.835 1.765 6.48 2.19 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.7001 ;
  ANTENNAPARTIALMETALAREA 0.5997 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.915 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.315 1.19 15.37 1.53 ;
      RECT 15.215 1.165 15.315 1.53 ;
      RECT 14.985 1.165 15.215 2.94 ;
      RECT 14.755 2.71 14.985 3.28 ;
      RECT 14.735 2.965 14.755 3.225 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.6464 ;
  ANTENNAPARTIALMETALAREA 0.9967 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9644 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.915 2.955 16.945 3.23 ;
      RECT 16.895 1.105 16.915 3.23 ;
      RECT 16.89 1.105 16.895 4.14 ;
      RECT 16.685 1.05 16.89 4.14 ;
      RECT 16.55 1.05 16.685 1.39 ;
      RECT 16.635 2.965 16.685 4.14 ;
      RECT 16.43 3.2 16.635 4.14 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.437 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4045 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.04 0.845 2.66 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1944 ;
  ANTENNAPARTIALMETALAREA 0.3843 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3144 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.215 2.045 1.84 2.66 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.13 -0.4 17.16 0.4 ;
      RECT 15.79 -0.4 16.13 1.69 ;
      RECT 14.395 -0.4 15.79 0.4 ;
      RECT 14.055 -0.4 14.395 0.575 ;
      RECT 11.355 -0.4 14.055 0.4 ;
      RECT 11.015 -0.4 11.355 0.575 ;
      RECT 8.785 -0.4 11.015 0.4 ;
      RECT 8.445 -0.4 8.785 1.37 ;
      RECT 7.01 -0.4 8.445 0.4 ;
      RECT 6.78 -0.4 7.01 0.9 ;
      RECT 4.095 -0.4 6.78 0.4 ;
      RECT 3.755 -0.4 4.095 0.9 ;
      RECT 1.18 -0.4 3.755 0.4 ;
      RECT 0.84 -0.4 1.18 0.575 ;
      RECT 0 -0.4 0.84 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.95 4.64 17.16 5.44 ;
      RECT 15.61 4.09 15.95 5.44 ;
      RECT 13.37 4.64 15.61 5.44 ;
      RECT 13.03 3.56 13.37 5.44 ;
      RECT 12.285 4.64 13.03 5.44 ;
      RECT 12.055 3.485 12.285 5.44 ;
      RECT 10.785 3.485 12.055 3.715 ;
      RECT 5.38 4.64 12.055 5.44 ;
      RECT 10.555 3.485 10.785 3.845 ;
      RECT 8.845 3.615 10.555 3.845 ;
      RECT 8.615 3.515 8.845 3.845 ;
      RECT 8.375 3.515 8.615 3.745 ;
      RECT 5.04 4.465 5.38 5.44 ;
      RECT 4.155 4.64 5.04 5.44 ;
      RECT 3.815 4.465 4.155 5.44 ;
      RECT 1.165 4.64 3.815 5.44 ;
      RECT 0.825 4.465 1.165 5.44 ;
      RECT 0 4.64 0.825 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.825 2.145 16.33 2.375 ;
      RECT 15.595 2.145 15.825 3.83 ;
      RECT 14.455 3.6 15.595 3.83 ;
      RECT 14.43 3.6 14.455 3.895 ;
      RECT 14.415 1.225 14.43 3.95 ;
      RECT 14.2 1.17 14.415 3.95 ;
      RECT 14.075 1.17 14.2 1.51 ;
      RECT 14.095 3.665 14.2 3.95 ;
      RECT 13.755 3.665 14.095 4.005 ;
      RECT 13.685 1.825 13.915 3.165 ;
      RECT 12.9 1.825 13.685 2.055 ;
      RECT 11.695 2.935 13.685 3.165 ;
      RECT 13.54 0.78 13.595 1.12 ;
      RECT 13.255 0.745 13.54 1.12 ;
      RECT 12.155 0.745 13.255 0.975 ;
      RECT 12.67 1.275 12.9 2.055 ;
      RECT 12.535 1.275 12.67 1.505 ;
      RECT 12.07 1.855 12.3 2.23 ;
      RECT 11.87 0.745 12.155 1.12 ;
      RECT 10.945 1.855 12.07 2.085 ;
      RECT 11.815 0.78 11.87 1.12 ;
      RECT 11.465 2.615 11.695 3.165 ;
      RECT 10.61 2.615 11.465 2.845 ;
      RECT 10.715 1.335 10.945 2.085 ;
      RECT 10.295 1.335 10.715 1.565 ;
      RECT 9.44 0.735 10.585 0.965 ;
      RECT 10.065 1.335 10.295 3.325 ;
      RECT 9.725 1.28 10.065 1.62 ;
      RECT 9.655 3.095 10.065 3.325 ;
      RECT 9.455 2.525 9.75 2.755 ;
      RECT 9.44 1.6 9.455 2.755 ;
      RECT 9.42 0.735 9.44 2.755 ;
      RECT 9.21 0.735 9.42 3.285 ;
      RECT 7.93 1.6 9.21 1.83 ;
      RECT 9.19 2.525 9.21 3.285 ;
      RECT 7.94 3.055 9.19 3.285 ;
      RECT 8.73 2.06 8.96 2.515 ;
      RECT 7.47 2.06 8.73 2.29 ;
      RECT 7.48 2.525 8.115 2.755 ;
      RECT 7.71 3.055 7.94 3.8 ;
      RECT 7.7 0.63 7.93 1.83 ;
      RECT 7.495 0.63 7.7 0.86 ;
      RECT 7.25 2.525 7.48 3.89 ;
      RECT 7.24 1.135 7.47 2.29 ;
      RECT 6.305 3.66 7.25 3.89 ;
      RECT 5.57 1.135 7.24 1.365 ;
      RECT 6.78 1.6 7.01 3.375 ;
      RECT 6.535 2.905 6.78 3.375 ;
      RECT 5.91 2.905 6.535 3.135 ;
      RECT 6.075 3.545 6.305 3.89 ;
      RECT 3.72 3.545 6.075 3.775 ;
      RECT 5.68 2.5 5.91 3.135 ;
      RECT 5.45 1.12 5.57 1.46 ;
      RECT 5.22 1.12 5.45 3.315 ;
      RECT 3.89 3.085 5.22 3.315 ;
      RECT 4.76 1.65 4.99 2.205 ;
      RECT 3.43 1.975 4.76 2.205 ;
      RECT 3.66 2.5 3.89 3.315 ;
      RECT 3.49 3.545 3.72 3.83 ;
      RECT 2.52 3.6 3.49 3.83 ;
      RECT 3.2 1.01 3.43 2.965 ;
      RECT 2.935 1.01 3.2 1.24 ;
      RECT 2.98 2.735 3.2 2.965 ;
      RECT 2.75 2.735 2.98 3.37 ;
      RECT 2.335 1.77 2.97 2.115 ;
      RECT 2.595 0.9 2.935 1.24 ;
      RECT 2.335 3.28 2.52 3.83 ;
      RECT 2.29 1.51 2.335 3.83 ;
      RECT 2.14 1.51 2.29 3.645 ;
      RECT 2.105 1.51 2.14 3.535 ;
      RECT 1.965 1.51 2.105 1.75 ;
      RECT 1.625 3.305 2.105 3.535 ;
      RECT 1.7 0.635 2.075 1.055 ;
      RECT 1.735 3.96 2.06 4.38 ;
      RECT 1.625 1.41 1.965 1.75 ;
      RECT 0.605 3.96 1.735 4.19 ;
      RECT 0.51 0.825 1.7 1.055 ;
      RECT 0.375 3.06 0.605 4.19 ;
      RECT 0.28 0.825 0.51 1.75 ;
      RECT 0.265 3.06 0.375 3.4 ;
  END
END DFFNSRX2

MACRO DFFNSRX1
  CLASS CORE ;
  FOREIGN DFFNSRX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 16.5 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSRXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3312 ;
  ANTENNAPARTIALMETALAREA 1.8312 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.5436 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.505 4.035 11.665 4.365 ;
      RECT 11.275 3.98 11.505 4.365 ;
      RECT 8.55 4.135 11.275 4.365 ;
      RECT 8.32 4.125 8.55 4.365 ;
      RECT 5.745 4.125 8.32 4.355 ;
      RECT 5.515 4.005 5.745 4.355 ;
      RECT 4.59 4.005 5.515 4.235 ;
      RECT 4.25 4.005 4.59 4.365 ;
     END
  END SN

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.3159 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.65 1.785 6.46 2.175 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6144 ;
  ANTENNAPARTIALMETALAREA 0.5568 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6606 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.595 2.94 14.965 3.225 ;
      RECT 14.595 1.46 14.65 1.8 ;
      RECT 14.365 1.46 14.595 3.225 ;
      RECT 14.31 1.46 14.365 1.8 ;
      RECT 14.33 2.995 14.365 3.225 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.84 ;
  ANTENNAPARTIALMETALAREA 0.777 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4927 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.21 2.94 16.285 3.705 ;
      RECT 16.07 1.48 16.21 3.705 ;
      RECT 15.98 1.48 16.07 3.76 ;
      RECT 15.97 1.48 15.98 1.71 ;
      RECT 15.73 3.42 15.98 3.76 ;
      RECT 15.63 1.37 15.97 1.71 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.3628 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4204 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 2.28 0.57 2.62 ;
      RECT 0.14 2.085 0.52 2.995 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.5415 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.59 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.38 1.695 2.985 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.21 -0.4 16.5 0.4 ;
      RECT 14.87 -0.4 15.21 0.575 ;
      RECT 11.27 -0.4 14.87 0.4 ;
      RECT 10.93 -0.4 11.27 0.575 ;
      RECT 8.705 -0.4 10.93 0.4 ;
      RECT 8.365 -0.4 8.705 1.38 ;
      RECT 6.755 -0.4 8.365 0.4 ;
      RECT 6.525 -0.4 6.755 0.9 ;
      RECT 3.96 -0.4 6.525 0.4 ;
      RECT 3.62 -0.4 3.96 0.9 ;
      RECT 1.23 -0.4 3.62 0.4 ;
      RECT 0.89 -0.4 1.23 0.575 ;
      RECT 0 -0.4 0.89 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.51 4.64 16.5 5.44 ;
      RECT 15.17 4.465 15.51 5.44 ;
      RECT 13.4 4.64 15.17 5.44 ;
      RECT 13.06 3.65 13.4 5.44 ;
      RECT 12.2 4.64 13.06 5.44 ;
      RECT 11.97 3.43 12.2 5.44 ;
      RECT 10.735 3.43 11.97 3.66 ;
      RECT 5.28 4.64 11.97 5.44 ;
      RECT 10.505 3.43 10.735 3.845 ;
      RECT 8.795 3.615 10.505 3.845 ;
      RECT 8.565 3.52 8.795 3.845 ;
      RECT 8.285 3.52 8.565 3.75 ;
      RECT 4.94 4.465 5.28 5.44 ;
      RECT 4.02 4.64 4.94 5.44 ;
      RECT 3.68 4.465 4.02 5.44 ;
      RECT 1.12 4.64 3.68 5.44 ;
      RECT 0.78 4.465 1.12 5.44 ;
      RECT 0 4.64 0.78 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.5 2.145 15.61 2.375 ;
      RECT 15.27 2.145 15.5 3.69 ;
      RECT 13.96 3.46 15.27 3.69 ;
      RECT 13.96 0.63 14.01 2.23 ;
      RECT 13.78 0.63 13.96 3.69 ;
      RECT 13.67 0.63 13.78 0.86 ;
      RECT 13.73 2 13.78 3.69 ;
      RECT 13.62 2.88 13.73 3.22 ;
      RECT 12.775 2.31 13.495 2.65 ;
      RECT 13.24 1.385 13.455 1.73 ;
      RECT 13.225 0.63 13.24 1.73 ;
      RECT 13.01 0.63 13.225 1.615 ;
      RECT 12.03 0.63 13.01 0.86 ;
      RECT 12.545 1.09 12.775 3.165 ;
      RECT 12.41 1.09 12.545 1.32 ;
      RECT 11.645 2.935 12.545 3.165 ;
      RECT 11.98 1.855 12.21 2.23 ;
      RECT 11.8 0.63 12.03 1.29 ;
      RECT 10.08 1.855 11.98 2.085 ;
      RECT 11.69 0.95 11.8 1.29 ;
      RECT 11.415 2.615 11.645 3.165 ;
      RECT 10.555 2.615 11.415 2.845 ;
      RECT 10.46 0.715 10.515 0.945 ;
      RECT 10.23 0.71 10.46 0.945 ;
      RECT 9.375 0.71 10.23 0.94 ;
      RECT 9.85 1.175 10.08 3.33 ;
      RECT 9.81 1.175 9.85 2.085 ;
      RECT 9.605 3.1 9.85 3.33 ;
      RECT 9.645 1.175 9.81 1.405 ;
      RECT 9.375 2.525 9.615 2.755 ;
      RECT 9.37 0.71 9.375 2.755 ;
      RECT 9.145 0.71 9.37 3.225 ;
      RECT 7.85 1.615 9.145 1.845 ;
      RECT 9.14 2.525 9.145 3.225 ;
      RECT 7.85 2.995 9.14 3.225 ;
      RECT 8.57 2.075 8.8 2.605 ;
      RECT 7.39 2.075 8.57 2.305 ;
      RECT 7.39 2.535 8.185 2.765 ;
      RECT 7.62 0.675 7.85 1.845 ;
      RECT 7.62 2.995 7.85 3.8 ;
      RECT 7.41 0.675 7.62 0.905 ;
      RECT 7.16 1.135 7.39 2.305 ;
      RECT 7.16 2.535 7.39 3.845 ;
      RECT 5.4 1.135 7.16 1.365 ;
      RECT 6.205 3.615 7.16 3.845 ;
      RECT 6.92 2.555 6.93 2.895 ;
      RECT 6.78 1.635 6.92 2.895 ;
      RECT 6.69 1.635 6.78 3.375 ;
      RECT 6.495 2.555 6.69 3.375 ;
      RECT 6.44 2.905 6.495 3.375 ;
      RECT 5.775 2.905 6.44 3.135 ;
      RECT 5.975 3.515 6.205 3.845 ;
      RECT 3.315 3.515 5.975 3.745 ;
      RECT 5.545 2.54 5.775 3.135 ;
      RECT 5.315 1.12 5.4 1.46 ;
      RECT 5.085 1.12 5.315 3.135 ;
      RECT 5.06 1.12 5.085 1.46 ;
      RECT 4.82 2.905 5.085 3.135 ;
      RECT 4.625 1.84 4.855 2.205 ;
      RECT 3.755 2.905 4.82 3.26 ;
      RECT 3.295 1.975 4.625 2.205 ;
      RECT 3.525 2.51 3.755 3.26 ;
      RECT 3.085 3.515 3.315 4.41 ;
      RECT 3.065 0.955 3.295 2.965 ;
      RECT 2.385 4.18 3.085 4.41 ;
      RECT 2.73 0.955 3.065 1.24 ;
      RECT 2.845 2.735 3.065 2.965 ;
      RECT 2.615 2.735 2.845 3.525 ;
      RECT 2.385 1.77 2.835 2.11 ;
      RECT 2.39 0.9 2.73 1.24 ;
      RECT 2.155 1.485 2.385 4.41 ;
      RECT 1.92 1.485 2.155 1.72 ;
      RECT 1.54 3.25 2.155 3.535 ;
      RECT 1.69 0.695 1.93 0.925 ;
      RECT 1.6 4.005 1.925 4.38 ;
      RECT 1.58 1.38 1.92 1.72 ;
      RECT 1.46 0.695 1.69 1.04 ;
      RECT 0.52 4.005 1.6 4.235 ;
      RECT 0.465 0.81 1.46 1.04 ;
      RECT 0.29 3.4 0.52 4.235 ;
      RECT 0.235 0.81 0.465 1.72 ;
      RECT 0.18 3.4 0.29 3.74 ;
  END
END DFFNSRX1

MACRO DFFNSXL
  CLASS CORE ;
  FOREIGN DFFNSXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.3192 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1978 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.115 3.77 10.675 4.34 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.53 ;
  ANTENNAPARTIALMETALAREA 1.2905 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.1056 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.655 0.865 12.885 3.755 ;
      RECT 12.255 0.865 12.655 1.095 ;
      RECT 12.395 3.5 12.655 3.755 ;
      RECT 12.325 3.525 12.395 3.755 ;
      RECT 12.095 3.525 12.325 3.85 ;
      RECT 12.025 0.745 12.255 1.095 ;
      RECT 12.07 3.62 12.095 3.85 ;
      RECT 11.84 3.62 12.07 4.195 ;
      RECT 11.5 0.745 12.025 0.975 ;
      RECT 11.73 3.855 11.84 4.195 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5172 ;
  ANTENNAPARTIALMETALAREA 0.8297 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0475 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.42 1.21 13.66 3.25 ;
      RECT 13.34 1.21 13.42 3.435 ;
      RECT 13.185 1.21 13.34 1.59 ;
      RECT 13.165 2.845 13.34 3.435 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2755 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.37 1.84 2.095 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2079 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9699 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.685 2.28 1.18 2.7 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.87 -0.4 13.86 0.4 ;
      RECT 12.53 -0.4 12.87 0.575 ;
      RECT 11.1 -0.4 12.53 0.4 ;
      RECT 10.76 -0.4 11.1 1.03 ;
      RECT 9.04 -0.4 10.76 0.4 ;
      RECT 8.7 -0.4 9.04 0.575 ;
      RECT 6.47 -0.4 8.7 0.4 ;
      RECT 6.24 -0.4 6.47 1.135 ;
      RECT 4.16 -0.4 6.24 0.4 ;
      RECT 3.82 -0.4 4.16 1.065 ;
      RECT 1.275 -0.4 3.82 0.4 ;
      RECT 0.935 -0.4 1.275 0.575 ;
      RECT 0 -0.4 0.935 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.93 4.64 13.86 5.44 ;
      RECT 12.495 4.465 12.93 5.44 ;
      RECT 11.235 4.64 12.495 5.44 ;
      RECT 11.005 3.265 11.235 5.44 ;
      RECT 9.68 4.64 11.005 5.44 ;
      RECT 9.34 4.14 9.68 5.44 ;
      RECT 7.09 4.64 9.34 5.44 ;
      RECT 6.86 3.765 7.09 5.44 ;
      RECT 5.695 4.64 6.86 5.44 ;
      RECT 5.355 4.11 5.695 5.44 ;
      RECT 4.405 4.64 5.355 5.44 ;
      RECT 4.065 4.465 4.405 5.44 ;
      RECT 1.47 4.64 4.065 5.44 ;
      RECT 1.13 4.465 1.47 5.44 ;
      RECT 0 4.64 1.13 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.155 1.6 12.185 2.375 ;
      RECT 11.955 1.6 12.155 3.19 ;
      RECT 11.88 1.6 11.955 1.83 ;
      RECT 11.925 2.075 11.955 3.19 ;
      RECT 11.71 2.96 11.925 3.19 ;
      RECT 11.54 1.49 11.88 1.83 ;
      RECT 11.11 2.14 11.45 2.48 ;
      RECT 10.515 2.195 11.11 2.425 ;
      RECT 10.49 1.62 10.515 3.375 ;
      RECT 10.285 1.62 10.49 3.43 ;
      RECT 9.74 1.62 10.285 1.85 ;
      RECT 10.15 3.09 10.285 3.43 ;
      RECT 8.5 2.435 10.03 2.665 ;
      RECT 9.4 1.19 9.74 1.85 ;
      RECT 9.21 1.62 9.4 1.85 ;
      RECT 8.87 1.62 9.21 1.96 ;
      RECT 8.465 1.545 8.5 3.835 ;
      RECT 8.27 1.545 8.465 3.89 ;
      RECT 7.215 0.675 8.29 0.905 ;
      RECT 7.825 1.545 8.27 1.775 ;
      RECT 8.125 3.55 8.27 3.89 ;
      RECT 7.215 2.515 8.04 2.915 ;
      RECT 7.595 1.19 7.825 1.775 ;
      RECT 6.985 0.675 7.215 2.915 ;
      RECT 6.01 1.37 6.985 1.6 ;
      RECT 6.445 2.685 6.985 2.915 ;
      RECT 5.795 1.855 6.755 2.085 ;
      RECT 6.215 2.685 6.445 3.405 ;
      RECT 5.945 3.65 6.175 4.04 ;
      RECT 5.78 0.695 6.01 1.6 ;
      RECT 3.61 3.65 5.945 3.88 ;
      RECT 5.565 1.855 5.795 3.415 ;
      RECT 4.71 0.63 5.78 0.925 ;
      RECT 5.55 1.855 5.565 2.085 ;
      RECT 4.465 3.185 5.565 3.415 ;
      RECT 5.32 1.45 5.55 2.085 ;
      RECT 5.095 2.355 5.325 2.74 ;
      RECT 4.985 2.355 5.095 2.585 ;
      RECT 4.755 1.32 4.985 2.585 ;
      RECT 3.575 1.32 4.755 1.55 ;
      RECT 4.655 0.63 4.71 0.86 ;
      RECT 4.235 2.035 4.465 3.415 ;
      RECT 3.755 2.035 4.235 2.265 ;
      RECT 3.38 2.57 3.61 4.205 ;
      RECT 3.345 1.13 3.575 1.55 ;
      RECT 3.305 2.57 3.38 2.8 ;
      RECT 1.96 3.975 3.38 4.205 ;
      RECT 2.795 1.13 3.345 1.36 ;
      RECT 3.105 1.885 3.305 2.8 ;
      RECT 2.895 3.035 3.125 3.52 ;
      RECT 3.075 1.6 3.105 2.8 ;
      RECT 2.82 1.6 3.075 2.115 ;
      RECT 2.84 3.035 2.895 3.265 ;
      RECT 2.61 2.595 2.84 3.265 ;
      RECT 2.505 0.87 2.795 1.36 ;
      RECT 2.505 2.595 2.61 2.825 ;
      RECT 2.455 0.87 2.505 2.825 ;
      RECT 2.275 1.13 2.455 2.825 ;
      RECT 1.73 3.945 1.96 4.205 ;
      RECT 0.395 3.945 1.73 4.175 ;
      RECT 0.395 1.195 0.54 1.535 ;
      RECT 0.395 3.295 0.52 3.635 ;
      RECT 0.2 1.195 0.395 4.175 ;
      RECT 0.165 1.225 0.2 4.175 ;
  END
END DFFNSXL

MACRO DFFNSX4
  CLASS CORE ;
  FOREIGN DFFNSX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 19.14 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9288 ;
  ANTENNAPARTIALMETALAREA 0.2356 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.47 4.01 5.09 4.39 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4225 ;
  ANTENNAPARTIALMETALAREA 0.9871 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2595 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.02 2.875 17.035 3.215 ;
      RECT 16.8 1.2 17.02 3.215 ;
      RECT 16.695 0.715 16.8 3.215 ;
      RECT 16.64 0.715 16.695 2.66 ;
      RECT 16.46 0.715 16.64 1.655 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4225 ;
  ANTENNAPARTIALMETALAREA 0.9892 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0846 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.34 0.955 18.35 2.7 ;
      RECT 18.24 0.955 18.34 3.22 ;
      RECT 17.96 0.76 18.24 3.22 ;
      RECT 17.955 0.76 17.96 3.16 ;
      RECT 17.9 0.76 17.955 1.57 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.162 ;
  ANTENNAPARTIALMETALAREA 0.2325 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.59 1.445 1.93 2.09 ;
      RECT 1.535 1.835 1.59 2.075 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.76 2.055 1.17 2.66 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.96 -0.4 19.14 0.4 ;
      RECT 18.62 -0.4 18.96 1.565 ;
      RECT 17.52 -0.4 18.62 0.4 ;
      RECT 17.18 -0.4 17.52 0.96 ;
      RECT 16.04 -0.4 17.18 0.4 ;
      RECT 15.7 -0.4 16.04 0.915 ;
      RECT 14.78 -0.4 15.7 0.4 ;
      RECT 14.44 -0.4 14.78 1.19 ;
      RECT 12.175 -0.4 14.44 0.4 ;
      RECT 11.835 -0.4 12.175 0.575 ;
      RECT 10.1 -0.4 11.835 0.4 ;
      RECT 9.76 -0.4 10.1 0.575 ;
      RECT 7.42 -0.4 9.76 0.4 ;
      RECT 7.08 -0.4 7.42 1.08 ;
      RECT 4.375 -0.4 7.08 0.4 ;
      RECT 4.035 -0.4 4.375 1.225 ;
      RECT 1.395 -0.4 4.035 0.4 ;
      RECT 1.055 -0.4 1.395 0.575 ;
      RECT 0 -0.4 1.055 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.955 4.64 19.14 5.44 ;
      RECT 18.615 4.055 18.955 5.44 ;
      RECT 17.675 4.64 18.615 5.44 ;
      RECT 17.335 4.015 17.675 5.44 ;
      RECT 16.395 4.64 17.335 5.44 ;
      RECT 16.055 4.055 16.395 5.44 ;
      RECT 14.97 4.64 16.055 5.44 ;
      RECT 14.63 3.52 14.97 5.44 ;
      RECT 13.53 4.64 14.63 5.44 ;
      RECT 13.19 3.52 13.53 5.44 ;
      RECT 12.05 4.64 13.19 5.44 ;
      RECT 11.71 4.015 12.05 5.44 ;
      RECT 9.98 4.64 11.71 5.44 ;
      RECT 9.64 3.38 9.98 5.44 ;
      RECT 7.38 4.64 9.64 5.44 ;
      RECT 7.04 3.33 7.38 5.44 ;
      RECT 5.72 4.64 7.04 5.44 ;
      RECT 5.38 4.195 5.72 5.44 ;
      RECT 4.175 4.64 5.38 5.44 ;
      RECT 3.945 4.15 4.175 5.44 ;
      RECT 1.39 4.64 3.945 5.44 ;
      RECT 1.05 4.465 1.39 5.44 ;
      RECT 0 4.64 1.05 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 18.645 2.06 18.875 3.725 ;
      RECT 16.115 3.495 18.645 3.725 ;
      RECT 15.885 1.62 16.115 3.725 ;
      RECT 15.5 1.62 15.885 1.85 ;
      RECT 15.69 3.055 15.885 3.725 ;
      RECT 15.35 3.055 15.69 3.865 ;
      RECT 15.215 1.28 15.5 1.85 ;
      RECT 14.25 2.08 15.46 2.42 ;
      RECT 15.16 1.28 15.215 1.62 ;
      RECT 14.195 2.08 14.25 3.34 ;
      RECT 14.02 1.505 14.195 3.34 ;
      RECT 13.965 1.505 14.02 2.31 ;
      RECT 13.91 2.975 14.02 3.34 ;
      RECT 13.59 1.505 13.965 1.735 ;
      RECT 12.81 2.975 13.91 3.205 ;
      RECT 13.28 2.13 13.62 2.47 ;
      RECT 13.525 1.295 13.59 1.735 ;
      RECT 13.36 1.055 13.525 1.735 ;
      RECT 13.16 1.055 13.36 1.58 ;
      RECT 10.855 2.185 13.28 2.415 ;
      RECT 11.435 1.055 13.16 1.285 ;
      RECT 12.7 2.975 12.81 3.34 ;
      RECT 12.47 2.975 12.7 3.725 ;
      RECT 11.46 3.495 12.47 3.725 ;
      RECT 11.23 3.495 11.46 4.04 ;
      RECT 9.405 0.865 10.975 1.095 ;
      RECT 10.63 1.385 10.855 3.085 ;
      RECT 10.625 1.385 10.63 3.26 ;
      RECT 10.355 1.385 10.625 1.77 ;
      RECT 10.4 2.855 10.625 3.26 ;
      RECT 8.66 2.915 10.4 3.145 ;
      RECT 10.08 2.275 10.39 2.505 ;
      RECT 8.94 1.385 10.355 1.615 ;
      RECT 9.85 2.175 10.08 2.505 ;
      RECT 9.505 2.175 9.85 2.405 ;
      RECT 9.275 1.925 9.505 2.405 ;
      RECT 9.175 0.675 9.405 1.095 ;
      RECT 8.74 1.925 9.275 2.155 ;
      RECT 8.1 0.675 9.175 0.905 ;
      RECT 8.71 1.195 8.94 1.615 ;
      RECT 8.4 1.195 8.71 1.425 ;
      RECT 8.375 2.915 8.66 3.44 ;
      RECT 8.015 2.31 8.41 2.65 ;
      RECT 8.32 3.1 8.375 3.44 ;
      RECT 8.015 0.675 8.1 1.625 ;
      RECT 7.87 0.675 8.015 3.1 ;
      RECT 7.785 1.395 7.87 3.1 ;
      RECT 6.62 1.395 7.785 1.645 ;
      RECT 6.705 2.87 7.785 3.1 ;
      RECT 6.215 2.235 7.495 2.635 ;
      RECT 6.475 2.87 6.705 3.265 ;
      RECT 6.335 0.675 6.62 1.645 ;
      RECT 6.105 3.035 6.475 3.265 ;
      RECT 6.115 3.52 6.345 4.1 ;
      RECT 6.28 0.675 6.335 1.6 ;
      RECT 6.18 0.675 6.28 1.04 ;
      RECT 5.815 2.23 6.215 2.635 ;
      RECT 3.515 3.52 6.115 3.75 ;
      RECT 5.71 1.715 5.815 3.265 ;
      RECT 5.585 1.015 5.71 3.265 ;
      RECT 5.48 1.015 5.585 1.945 ;
      RECT 4.09 3.035 5.585 3.265 ;
      RECT 5.315 1.015 5.48 1.245 ;
      RECT 5.005 2.455 5.29 2.685 ;
      RECT 4.775 1.495 5.005 2.685 ;
      RECT 3.015 1.495 4.775 1.725 ;
      RECT 3.86 2.01 4.09 3.265 ;
      RECT 3.285 2.075 3.515 4.345 ;
      RECT 3.065 2.075 3.285 2.305 ;
      RECT 1.885 4.115 3.285 4.345 ;
      RECT 2.835 3 3.05 3.71 ;
      RECT 2.905 1 3.015 1.725 ;
      RECT 2.835 1 2.905 1.84 ;
      RECT 2.82 1 2.835 3.71 ;
      RECT 2.675 1 2.82 3.23 ;
      RECT 2.605 1.61 2.675 3.23 ;
      RECT 1.655 3.875 1.885 4.345 ;
      RECT 0.465 3.875 1.655 4.105 ;
      RECT 0.465 1.27 0.52 1.61 ;
      RECT 0.465 2.96 0.52 3.3 ;
      RECT 0.235 1.27 0.465 4.105 ;
      RECT 0.18 1.27 0.235 1.61 ;
      RECT 0.18 2.96 0.235 3.3 ;
  END
END DFFNSX4

MACRO DFFNSX2
  CLASS CORE ;
  FOREIGN DFFNSX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.522 ;
  ANTENNAPARTIALMETALAREA 0.2935 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.76 3.95 10.405 4.405 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.088 ;
  ANTENNAPARTIALMETALAREA 0.647 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2065 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.145 0.835 12.325 2.92 ;
      RECT 12.13 0.69 12.145 2.92 ;
      RECT 12.095 0.69 12.13 3.11 ;
      RECT 11.915 0.69 12.095 1.065 ;
      RECT 12.02 2.635 12.095 3.11 ;
      RECT 11.9 2.69 12.02 3.11 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4592 ;
  ANTENNAPARTIALMETALAREA 0.9442 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.293 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.645 1.845 13.72 3.13 ;
      RECT 13.64 0.955 13.645 3.13 ;
      RECT 13.575 0.755 13.64 3.13 ;
      RECT 13.49 0.755 13.575 4.24 ;
      RECT 13.415 0.755 13.49 2.075 ;
      RECT 13.345 2.9 13.49 4.24 ;
      RECT 13.3 0.755 13.415 1.565 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3309 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2879 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.38 1.84 1.97 ;
      RECT 1.535 1.38 1.765 2.075 ;
      RECT 1.32 1.38 1.535 1.97 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.2704 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.66 2.32 1.18 2.84 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.92 -0.4 13.86 0.4 ;
      RECT 12.58 -0.4 12.92 1.475 ;
      RECT 11.06 -0.4 12.58 0.4 ;
      RECT 10.72 -0.4 11.06 0.575 ;
      RECT 9.04 -0.4 10.72 0.4 ;
      RECT 8.7 -0.4 9.04 0.575 ;
      RECT 6.47 -0.4 8.7 0.4 ;
      RECT 6.24 -0.4 6.47 1.135 ;
      RECT 4.16 -0.4 6.24 0.4 ;
      RECT 3.82 -0.4 4.16 1.065 ;
      RECT 1.4 -0.4 3.82 0.4 ;
      RECT 1.06 -0.4 1.4 0.575 ;
      RECT 0 -0.4 1.06 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.91 4.64 13.86 5.44 ;
      RECT 12.57 3.925 12.91 5.44 ;
      RECT 10.895 4.64 12.57 5.44 ;
      RECT 10.865 3.505 10.895 5.44 ;
      RECT 10.665 3.34 10.865 5.44 ;
      RECT 10.635 3.34 10.665 3.735 ;
      RECT 9.44 4.64 10.665 5.44 ;
      RECT 9.1 4.14 9.44 5.44 ;
      RECT 6.945 4.64 9.1 5.44 ;
      RECT 6.715 3.77 6.945 5.44 ;
      RECT 5.695 4.64 6.715 5.44 ;
      RECT 5.355 4.095 5.695 5.44 ;
      RECT 4.405 4.64 5.355 5.44 ;
      RECT 4.065 4.465 4.405 5.44 ;
      RECT 1.44 4.64 4.065 5.44 ;
      RECT 1.1 4.465 1.44 5.44 ;
      RECT 0 4.64 1.1 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.11 2.24 13.15 2.62 ;
      RECT 12.92 2.24 13.11 3.585 ;
      RECT 12.88 2.295 12.92 3.585 ;
      RECT 11.615 3.355 12.88 3.585 ;
      RECT 11.615 1.435 11.655 1.775 ;
      RECT 11.59 1.435 11.615 3.585 ;
      RECT 11.385 1.435 11.59 3.83 ;
      RECT 11.315 1.435 11.385 1.775 ;
      RECT 11.36 3.355 11.385 3.83 ;
      RECT 10.38 2.12 11.155 2.505 ;
      RECT 10.2 1.62 10.38 3.125 ;
      RECT 10.15 1.62 10.2 3.635 ;
      RECT 9.74 1.62 10.15 1.85 ;
      RECT 9.86 2.825 10.15 3.635 ;
      RECT 8.315 2.195 9.92 2.425 ;
      RECT 9.4 1.16 9.74 1.85 ;
      RECT 9.01 1.62 9.4 1.85 ;
      RECT 8.67 1.62 9.01 1.96 ;
      RECT 8.28 1.545 8.315 3.835 ;
      RECT 7.215 0.675 8.29 0.905 ;
      RECT 8.085 1.545 8.28 3.89 ;
      RECT 7.825 1.545 8.085 1.775 ;
      RECT 7.94 3.55 8.085 3.89 ;
      RECT 7.215 2.515 7.855 2.915 ;
      RECT 7.595 1.19 7.825 1.775 ;
      RECT 6.985 0.675 7.215 2.915 ;
      RECT 6.01 1.37 6.985 1.6 ;
      RECT 6.405 2.685 6.985 2.915 ;
      RECT 6.515 1.885 6.745 2.295 ;
      RECT 5.795 1.885 6.515 2.115 ;
      RECT 6.175 2.685 6.405 3.405 ;
      RECT 5.945 3.635 6.175 4.04 ;
      RECT 5.78 0.695 6.01 1.6 ;
      RECT 3.61 3.635 5.945 3.865 ;
      RECT 5.565 1.885 5.795 3.37 ;
      RECT 5.08 0.695 5.78 0.925 ;
      RECT 5.55 1.885 5.565 2.115 ;
      RECT 4.465 3.14 5.565 3.37 ;
      RECT 5.32 1.45 5.55 2.115 ;
      RECT 5.095 2.37 5.325 2.79 ;
      RECT 4.985 2.37 5.095 2.6 ;
      RECT 4.655 0.63 5.08 0.925 ;
      RECT 4.755 1.295 4.985 2.6 ;
      RECT 2.795 1.295 4.755 1.525 ;
      RECT 4.235 2.035 4.465 3.37 ;
      RECT 3.755 2.035 4.235 2.265 ;
      RECT 3.38 2.57 3.61 4.085 ;
      RECT 3.305 2.57 3.38 2.8 ;
      RECT 0.54 3.855 3.38 4.085 ;
      RECT 3.075 1.805 3.305 2.8 ;
      RECT 2.895 3.035 3.125 3.52 ;
      RECT 2.82 1.805 3.075 2.035 ;
      RECT 2.84 3.035 2.895 3.265 ;
      RECT 2.61 2.595 2.84 3.265 ;
      RECT 2.505 0.86 2.795 1.525 ;
      RECT 2.505 2.595 2.61 2.825 ;
      RECT 2.455 0.86 2.505 2.825 ;
      RECT 2.275 1.295 2.455 2.825 ;
      RECT 0.43 0.815 0.54 1.155 ;
      RECT 0.43 3.4 0.54 4.085 ;
      RECT 0.2 0.815 0.43 4.085 ;
  END
END DFFNSX2

MACRO DFFNSX1
  CLASS CORE ;
  FOREIGN DFFNSX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNSXL ;

  PIN SN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3348 ;
  ANTENNAPARTIALMETALAREA 0.3192 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1978 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.115 3.77 10.675 4.34 ;
     END
  END SN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.75 ;
  ANTENNAPARTIALMETALAREA 1.2699 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.0155 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.615 0.865 12.845 3.755 ;
      RECT 12.215 0.865 12.615 1.095 ;
      RECT 12.395 3.5 12.615 3.755 ;
      RECT 12.325 3.525 12.395 3.755 ;
      RECT 12.095 3.525 12.325 3.85 ;
      RECT 11.985 0.79 12.215 1.095 ;
      RECT 12.07 3.62 12.095 3.85 ;
      RECT 11.84 3.62 12.07 4.195 ;
      RECT 11.46 0.79 11.985 1.02 ;
      RECT 11.73 3.855 11.84 4.195 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.846 ;
  ANTENNAPARTIALMETALAREA 0.8711 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2754 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.415 1.21 13.66 3.25 ;
      RECT 13.34 1.21 13.415 3.67 ;
      RECT 13.185 1.21 13.34 1.59 ;
      RECT 13.185 2.845 13.34 3.67 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2755 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.375 1.84 2.1 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.18 ;
  ANTENNAPARTIALMETALAREA 0.2079 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9699 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.685 2.28 1.18 2.7 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.87 -0.4 13.86 0.4 ;
      RECT 12.53 -0.4 12.87 0.575 ;
      RECT 11.06 -0.4 12.53 0.4 ;
      RECT 10.72 -0.4 11.06 1.01 ;
      RECT 9.04 -0.4 10.72 0.4 ;
      RECT 8.7 -0.4 9.04 0.575 ;
      RECT 6.46 -0.4 8.7 0.4 ;
      RECT 6.23 -0.4 6.46 1.135 ;
      RECT 4.16 -0.4 6.23 0.4 ;
      RECT 3.82 -0.4 4.16 1.065 ;
      RECT 1.24 -0.4 3.82 0.4 ;
      RECT 0.9 -0.4 1.24 0.575 ;
      RECT 0 -0.4 0.9 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.93 4.64 13.86 5.44 ;
      RECT 12.495 4.465 12.93 5.44 ;
      RECT 11.235 4.64 12.495 5.44 ;
      RECT 11.005 3.03 11.235 5.44 ;
      RECT 9.68 4.64 11.005 5.44 ;
      RECT 9.34 4.14 9.68 5.44 ;
      RECT 7.09 4.64 9.34 5.44 ;
      RECT 6.86 3.765 7.09 5.44 ;
      RECT 5.695 4.64 6.86 5.44 ;
      RECT 5.355 4.095 5.695 5.44 ;
      RECT 4.405 4.64 5.355 5.44 ;
      RECT 4.065 4.465 4.405 5.44 ;
      RECT 1.56 4.64 4.065 5.44 ;
      RECT 1.22 4.465 1.56 5.44 ;
      RECT 0 4.64 1.22 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.155 2.02 12.185 2.375 ;
      RECT 11.925 1.6 12.155 3.095 ;
      RECT 11.84 1.6 11.925 1.83 ;
      RECT 11.71 2.865 11.925 3.095 ;
      RECT 11.5 1.49 11.84 1.83 ;
      RECT 11.11 2.14 11.45 2.48 ;
      RECT 10.515 2.195 11.11 2.425 ;
      RECT 10.49 1.62 10.515 3.345 ;
      RECT 10.285 1.62 10.49 3.4 ;
      RECT 9.74 1.62 10.285 1.85 ;
      RECT 10.15 3.06 10.285 3.4 ;
      RECT 8.5 2.435 10.03 2.665 ;
      RECT 9.4 1.19 9.74 1.85 ;
      RECT 9.21 1.62 9.4 1.85 ;
      RECT 8.87 1.62 9.21 1.96 ;
      RECT 8.465 1.545 8.5 3.835 ;
      RECT 8.27 1.545 8.465 3.89 ;
      RECT 7.215 0.675 8.29 0.905 ;
      RECT 7.825 1.545 8.27 1.775 ;
      RECT 8.125 3.55 8.27 3.89 ;
      RECT 7.215 2.515 8.04 2.915 ;
      RECT 7.595 1.19 7.825 1.775 ;
      RECT 6.985 0.675 7.215 2.915 ;
      RECT 6 1.37 6.985 1.6 ;
      RECT 6.445 2.685 6.985 2.915 ;
      RECT 5.795 1.835 6.745 2.065 ;
      RECT 6.215 2.685 6.445 3.405 ;
      RECT 5.945 3.635 6.175 4.04 ;
      RECT 5.78 0.695 6 1.6 ;
      RECT 3.61 3.635 5.945 3.865 ;
      RECT 5.565 1.835 5.795 3.37 ;
      RECT 5.77 0.675 5.78 1.6 ;
      RECT 4.71 0.675 5.77 0.925 ;
      RECT 5.54 1.835 5.565 2.065 ;
      RECT 4.465 3.14 5.565 3.37 ;
      RECT 5.31 1.42 5.54 2.065 ;
      RECT 5.095 2.355 5.325 2.74 ;
      RECT 4.985 2.355 5.095 2.585 ;
      RECT 4.755 1.295 4.985 2.585 ;
      RECT 2.795 1.295 4.755 1.525 ;
      RECT 4.655 0.675 4.71 0.905 ;
      RECT 4.235 2.005 4.465 3.37 ;
      RECT 3.705 2.005 4.235 2.235 ;
      RECT 3.38 2.57 3.61 4.085 ;
      RECT 3.305 2.57 3.38 2.8 ;
      RECT 1.575 3.855 3.38 4.085 ;
      RECT 3.075 1.805 3.305 2.8 ;
      RECT 2.895 3.035 3.125 3.52 ;
      RECT 2.82 1.805 3.075 2.035 ;
      RECT 2.84 3.035 2.895 3.265 ;
      RECT 2.61 2.595 2.84 3.265 ;
      RECT 2.505 0.86 2.795 1.525 ;
      RECT 2.505 2.595 2.61 2.825 ;
      RECT 2.455 0.86 2.505 2.825 ;
      RECT 2.275 1.295 2.455 2.825 ;
      RECT 1.345 3.855 1.575 4.175 ;
      RECT 0.395 3.945 1.345 4.175 ;
      RECT 0.395 1.195 0.54 1.535 ;
      RECT 0.395 3.36 0.52 3.7 ;
      RECT 0.2 1.195 0.395 4.175 ;
      RECT 0.165 1.225 0.2 4.175 ;
  END
END DFFNSX1

MACRO DFFNRXL
  CLASS CORE ;
  FOREIGN DFFNRXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3783 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.7914 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.59 2.9 4.93 3.24 ;
      RECT 4.48 2.9 4.59 3.185 ;
      RECT 4.25 2.36 4.48 3.185 ;
      RECT 4.12 2.36 4.25 2.68 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5343 ;
  ANTENNAPARTIALMETALAREA 1.2354 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4855 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.125 0.865 14.355 4.035 ;
      RECT 13.77 0.865 14.125 1.095 ;
      RECT 13.975 3.5 14.125 4.035 ;
      RECT 13.85 3.805 13.975 4.035 ;
      RECT 13.51 3.805 13.85 4.23 ;
      RECT 13.43 0.635 13.77 1.095 ;
      RECT 13.47 3.805 13.51 4.175 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 1.0166 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9379 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.495 3.62 15.58 3.96 ;
      RECT 15.265 1.89 15.495 3.96 ;
      RECT 15.18 1.89 15.265 2.12 ;
      RECT 15.24 3.62 15.265 3.96 ;
      RECT 14.66 1.19 15.18 2.12 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2509 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.525 1.575 1.915 2.105 ;
      RECT 1.455 1.715 1.525 2.08 ;
      RECT 1.4 1.74 1.455 2.08 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.5514 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.1147 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.91 2.635 1.23 3.22 ;
      RECT 0.91 1.885 1.02 2.405 ;
      RECT 0.68 1.885 0.91 3.22 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.5 -0.4 15.84 0.4 ;
      RECT 14.16 -0.4 14.5 0.575 ;
      RECT 12.89 -0.4 14.16 0.4 ;
      RECT 12.55 -0.4 12.89 0.95 ;
      RECT 11.13 -0.4 12.55 0.4 ;
      RECT 10.79 -0.4 11.13 1.11 ;
      RECT 6.365 -0.4 10.79 0.4 ;
      RECT 7.895 1.205 8.235 1.76 ;
      RECT 6.66 1.205 7.895 1.435 ;
      RECT 6.365 1.205 6.66 1.58 ;
      RECT 6.32 -0.4 6.365 1.58 ;
      RECT 6.135 -0.4 6.32 1.525 ;
      RECT 4.35 -0.4 6.135 0.4 ;
      RECT 4.01 -0.4 4.35 0.96 ;
      RECT 1.35 -0.4 4.01 0.4 ;
      RECT 1.01 -0.4 1.35 0.575 ;
      RECT 0 -0.4 1.01 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.81 4.64 15.84 5.44 ;
      RECT 14.47 4.465 14.81 5.44 ;
      RECT 13.09 4.64 14.47 5.44 ;
      RECT 12.75 4.11 13.09 5.44 ;
      RECT 11.065 4.64 12.75 5.44 ;
      RECT 10.725 4.08 11.065 5.44 ;
      RECT 8.73 4.64 10.725 5.44 ;
      RECT 7.79 4.08 8.73 5.44 ;
      RECT 4.66 4.64 7.79 5.44 ;
      RECT 4.32 4.465 4.66 5.44 ;
      RECT 1.65 4.64 4.32 5.44 ;
      RECT 1.31 4.08 1.65 5.44 ;
      RECT 0 4.64 1.31 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.74 1.38 13.85 3.16 ;
      RECT 13.51 1.38 13.74 3.35 ;
      RECT 13.33 1.38 13.51 1.85 ;
      RECT 13.4 2.82 13.51 3.35 ;
      RECT 12.985 1.88 13.03 2.22 ;
      RECT 12.975 1.865 12.985 2.22 ;
      RECT 12.475 1.865 12.975 2.245 ;
      RECT 12.245 1.865 12.475 3.85 ;
      RECT 12.035 1.865 12.245 2.095 ;
      RECT 11.77 3.62 12.245 3.85 ;
      RECT 11.805 0.915 12.035 2.095 ;
      RECT 11.67 3.005 12.01 3.39 ;
      RECT 11.645 0.915 11.805 1.825 ;
      RECT 11.43 3.62 11.77 3.96 ;
      RECT 10.535 3.16 11.67 3.39 ;
      RECT 11.235 1.595 11.645 1.825 ;
      RECT 11.235 2.24 11.29 2.58 ;
      RECT 11.005 1.595 11.235 2.58 ;
      RECT 10.95 2.24 11.005 2.58 ;
      RECT 10.355 1.425 10.535 3.405 ;
      RECT 10.355 4 10.36 4.34 ;
      RECT 10.305 1.425 10.355 4.34 ;
      RECT 9.59 1.425 10.305 1.655 ;
      RECT 10.125 3.16 10.305 4.34 ;
      RECT 10.02 4 10.125 4.34 ;
      RECT 9.615 2.39 9.955 2.73 ;
      RECT 9.53 0.63 9.87 0.97 ;
      RECT 8.935 2.445 9.615 2.675 ;
      RECT 9.305 1.29 9.59 1.655 ;
      RECT 8.935 0.685 9.53 0.915 ;
      RECT 9.25 1.29 9.305 1.63 ;
      RECT 8.705 0.675 8.935 3.465 ;
      RECT 7.315 0.675 8.705 0.915 ;
      RECT 8.15 3.075 8.705 3.465 ;
      RECT 6.975 2.14 8.39 2.48 ;
      RECT 7.855 2.81 7.91 3.15 ;
      RECT 7.625 2.81 7.855 3.825 ;
      RECT 7.57 2.81 7.625 3.15 ;
      RECT 7.495 3.595 7.625 3.825 ;
      RECT 7.265 3.595 7.495 4.365 ;
      RECT 7.03 0.675 7.315 0.905 ;
      RECT 5.125 4.135 7.265 4.365 ;
      RECT 6.69 0.635 7.03 0.975 ;
      RECT 6.745 1.825 6.975 3.69 ;
      RECT 5.71 1.825 6.745 2.055 ;
      RECT 6.44 3.46 6.745 3.69 ;
      RECT 6.1 3.46 6.44 3.8 ;
      RECT 6.09 2.44 6.43 2.78 ;
      RECT 5.485 2.495 6.09 2.725 ;
      RECT 5.71 1.1 5.72 1.44 ;
      RECT 5.48 1.1 5.71 2.055 ;
      RECT 5.485 3.485 5.705 3.87 ;
      RECT 5.365 2.435 5.485 3.87 ;
      RECT 5.38 1.1 5.48 1.885 ;
      RECT 3.9 1.655 5.38 1.885 ;
      RECT 5.255 2.435 5.365 3.715 ;
      RECT 5.25 2.435 5.255 2.665 ;
      RECT 4.915 2.115 5.25 2.665 ;
      RECT 4.895 3.945 5.125 4.365 ;
      RECT 4.895 0.77 5.12 1.11 ;
      RECT 4.91 2.115 4.915 2.455 ;
      RECT 4.78 0.77 4.895 1.42 ;
      RECT 4.005 3.945 4.895 4.175 ;
      RECT 4.665 0.825 4.78 1.42 ;
      RECT 2.86 1.19 4.665 1.42 ;
      RECT 3.795 2.935 4.005 4.355 ;
      RECT 3.56 1.655 3.9 2.055 ;
      RECT 3.775 2.395 3.795 4.355 ;
      RECT 3.565 2.395 3.775 3.165 ;
      RECT 2.93 4.125 3.775 4.355 ;
      RECT 3.235 2.395 3.565 2.625 ;
      RECT 3.535 1.655 3.56 2 ;
      RECT 3.275 3.46 3.46 3.8 ;
      RECT 3.045 2.935 3.275 3.8 ;
      RECT 3.005 1.705 3.235 2.625 ;
      RECT 2.695 2.935 3.045 3.165 ;
      RECT 2.895 1.705 3.005 2.055 ;
      RECT 2.59 4.07 2.93 4.41 ;
      RECT 2.84 1.715 2.895 2.055 ;
      RECT 2.525 0.9 2.86 1.42 ;
      RECT 2.525 2.545 2.695 3.165 ;
      RECT 2.385 4.07 2.59 4.355 ;
      RECT 2.465 0.9 2.525 3.165 ;
      RECT 2.295 0.9 2.465 2.775 ;
      RECT 2.155 3.62 2.385 4.355 ;
      RECT 0.6 3.62 2.155 3.85 ;
      RECT 0.45 3.51 0.6 3.85 ;
      RECT 0.45 1.04 0.56 1.38 ;
      RECT 0.22 1.04 0.45 3.85 ;
  END
END DFFNRXL

MACRO DFFNRX4
  CLASS CORE ;
  FOREIGN DFFNRX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.46 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4068 ;
  ANTENNAPARTIALMETALAREA 0.345 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.68 2.745 5.14 3.495 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2718 ;
  ANTENNAPARTIALMETALAREA 0.7831 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5917 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.96 1.195 18.34 3.22 ;
      RECT 17.94 1.195 17.96 1.535 ;
      RECT 17.94 2.78 17.96 3.12 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2718 ;
  ANTENNAPARTIALMETALAREA 0.7685 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5705 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 19.56 1.26 19.66 3.12 ;
      RECT 19.28 1.195 19.56 3.12 ;
      RECT 19.275 1.195 19.28 2.075 ;
      RECT 19.22 2.78 19.28 3.12 ;
      RECT 19.22 1.195 19.275 1.535 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.198 ;
  ANTENNAPARTIALMETALAREA 0.4378 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.6218 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.845 2.56 1.91 2.9 ;
      RECT 1.46 1.82 1.845 2.9 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2844 ;
  ANTENNAPARTIALMETALAREA 0.2886 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1395 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.66 2.175 1.18 2.73 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.2 -0.4 20.46 0.4 ;
      RECT 19.86 -0.4 20.2 0.95 ;
      RECT 18.92 -0.4 19.86 0.4 ;
      RECT 18.58 -0.4 18.92 0.95 ;
      RECT 17.64 -0.4 18.58 0.4 ;
      RECT 17.3 -0.4 17.64 0.95 ;
      RECT 16.27 -0.4 17.3 0.4 ;
      RECT 15.93 -0.4 16.27 0.95 ;
      RECT 14.83 -0.4 15.93 0.4 ;
      RECT 14.49 -0.4 14.83 0.95 ;
      RECT 13.37 -0.4 14.49 0.4 ;
      RECT 13.03 -0.4 13.37 0.95 ;
      RECT 11.6 -0.4 13.03 0.4 ;
      RECT 11.26 -0.4 11.6 0.575 ;
      RECT 9.005 -0.4 11.26 0.4 ;
      RECT 8.775 -0.4 9.005 1.475 ;
      RECT 7.15 -0.4 8.775 0.4 ;
      RECT 8.59 1.245 8.775 1.475 ;
      RECT 6.81 -0.4 7.15 0.96 ;
      RECT 5.14 -0.4 6.81 0.4 ;
      RECT 4.8 -0.4 5.14 1.335 ;
      RECT 1.08 -0.4 4.8 0.4 ;
      RECT 0.74 -0.4 1.08 0.575 ;
      RECT 0 -0.4 0.74 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.2 4.64 20.46 5.44 ;
      RECT 19.86 4.04 20.2 5.44 ;
      RECT 18.92 4.64 19.86 5.44 ;
      RECT 18.58 4.04 18.92 5.44 ;
      RECT 17.64 4.64 18.58 5.44 ;
      RECT 17.3 4.04 17.64 5.44 ;
      RECT 16.07 4.64 17.3 5.44 ;
      RECT 15.73 3.055 16.07 5.44 ;
      RECT 13.47 4.64 15.73 5.44 ;
      RECT 13.13 4.08 13.47 5.44 ;
      RECT 10.99 4.64 13.13 5.44 ;
      RECT 10.65 3.675 10.99 5.44 ;
      RECT 8.14 4.64 10.65 5.44 ;
      RECT 7.8 3.92 8.14 5.44 ;
      RECT 4.48 4.64 7.8 5.44 ;
      RECT 4.14 4.465 4.48 5.44 ;
      RECT 1.545 4.64 4.14 5.44 ;
      RECT 1.205 4.465 1.545 5.44 ;
      RECT 0 4.64 1.205 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 19.965 2.03 20.195 3.75 ;
      RECT 17.635 3.52 19.965 3.75 ;
      RECT 17.405 1.395 17.635 3.75 ;
      RECT 16.95 1.395 17.405 1.73 ;
      RECT 16.79 3.265 17.405 3.495 ;
      RECT 16.17 2.1 17.11 2.44 ;
      RECT 16.61 1.39 16.95 1.73 ;
      RECT 16.45 2.975 16.79 3.785 ;
      RECT 16.6 1.395 16.61 1.675 ;
      RECT 15.55 2.155 16.17 2.385 ;
      RECT 15.32 0.72 15.55 2.69 ;
      RECT 15.21 0.72 15.32 1.475 ;
      RECT 14.79 2.46 15.32 2.69 ;
      RECT 14.11 1.245 15.21 1.475 ;
      RECT 14.715 1.725 15.07 2.065 ;
      RECT 14.56 2.46 14.79 3.835 ;
      RECT 14.13 1.725 14.715 2.105 ;
      RECT 14.45 2.985 14.56 3.835 ;
      RECT 12.86 3.605 14.45 3.835 ;
      RECT 13.125 1.875 14.13 2.105 ;
      RECT 13.88 0.7 14.11 1.475 ;
      RECT 13.77 0.7 13.88 1.04 ;
      RECT 12.895 1.495 13.125 3.365 ;
      RECT 10.555 1.495 12.895 1.735 ;
      RECT 12.265 3.135 12.895 3.365 ;
      RECT 12.63 3.605 12.86 4.25 ;
      RECT 12.125 2.425 12.465 2.82 ;
      RECT 11.02 0.955 12.38 1.185 ;
      RECT 12.265 3.75 12.32 4.09 ;
      RECT 12.035 3.135 12.265 4.09 ;
      RECT 10.095 2.425 12.125 2.655 ;
      RECT 10.355 3.135 12.035 3.365 ;
      RECT 11.98 3.75 12.035 4.09 ;
      RECT 10.79 0.635 11.02 1.185 ;
      RECT 9.555 0.635 10.79 0.865 ;
      RECT 10.325 1.095 10.555 1.735 ;
      RECT 10.125 3.135 10.355 3.855 ;
      RECT 9.91 1.095 10.325 1.325 ;
      RECT 9.71 3.625 10.125 3.855 ;
      RECT 9.865 1.72 10.095 2.655 ;
      RECT 9.37 3.625 9.71 3.99 ;
      RECT 9.555 1.745 9.58 3.145 ;
      RECT 9.35 0.635 9.555 3.145 ;
      RECT 9.325 0.635 9.35 1.975 ;
      RECT 9.065 2.915 9.35 3.145 ;
      RECT 8.125 1.715 9.325 1.975 ;
      RECT 7.535 2.205 9.12 2.435 ;
      RECT 8.9 2.915 9.065 3.945 ;
      RECT 8.675 2.915 8.9 4 ;
      RECT 8.56 3.66 8.675 4 ;
      RECT 8.165 2.84 8.33 3.18 ;
      RECT 7.935 2.84 8.165 3.66 ;
      RECT 7.895 0.675 8.125 1.975 ;
      RECT 7.405 3.43 7.935 3.66 ;
      RECT 7.4 0.675 7.895 0.905 ;
      RECT 7.305 1.565 7.535 3.145 ;
      RECT 7.175 3.43 7.405 4.365 ;
      RECT 6.59 1.565 7.305 1.795 ;
      RECT 6.86 2.915 7.305 3.145 ;
      RECT 5.025 4.135 7.175 4.365 ;
      RECT 6.52 2.915 6.86 3.87 ;
      RECT 6.49 2.1 6.83 2.44 ;
      RECT 6.25 1.43 6.59 1.795 ;
      RECT 5.675 2.155 6.49 2.385 ;
      RECT 4.12 1.565 6.25 1.795 ;
      RECT 5.675 3.56 5.73 3.9 ;
      RECT 5.445 2.025 5.675 3.9 ;
      RECT 4.93 2.025 5.445 2.255 ;
      RECT 5.39 3.56 5.445 3.9 ;
      RECT 4.795 3.945 5.025 4.365 ;
      RECT 3.825 3.945 4.795 4.175 ;
      RECT 4.265 2.32 4.32 2.66 ;
      RECT 2.985 0.825 4.31 1.055 ;
      RECT 4.12 2.245 4.265 2.66 ;
      RECT 3.98 1.565 4.12 2.66 ;
      RECT 3.89 1.565 3.98 2.475 ;
      RECT 3.595 3.035 3.825 4.345 ;
      RECT 3.48 3.035 3.595 3.265 ;
      RECT 2.435 4.115 3.595 4.345 ;
      RECT 3.25 1.98 3.48 3.265 ;
      RECT 3.2 1.98 3.25 2.21 ;
      RECT 2.915 1.82 3.2 2.21 ;
      RECT 3.02 3.5 3.155 3.84 ;
      RECT 2.79 2.465 3.02 3.84 ;
      RECT 2.76 0.825 2.985 1.415 ;
      RECT 2.86 1.82 2.915 2.16 ;
      RECT 2.425 2.465 2.79 2.695 ;
      RECT 2.755 0.825 2.76 1.47 ;
      RECT 2.425 1.13 2.755 1.47 ;
      RECT 2.205 4.005 2.435 4.345 ;
      RECT 2.42 1.13 2.425 2.695 ;
      RECT 2.195 1.185 2.42 2.695 ;
      RECT 0.405 4.005 2.205 4.235 ;
      RECT 0.465 1.22 0.52 1.56 ;
      RECT 0.405 3.18 0.52 3.52 ;
      RECT 0.405 1.215 0.465 1.56 ;
      RECT 0.175 1.215 0.405 4.235 ;
  END
END DFFNRX4

MACRO DFFNRX2
  CLASS CORE ;
  FOREIGN DFFNRX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.3098 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.605 2.875 4.66 3.39 ;
      RECT 4.32 2.755 4.605 3.39 ;
      RECT 4.175 2.755 4.32 3.335 ;
      RECT 4.13 2.875 4.175 3.24 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1736 ;
  ANTENNAPARTIALMETALAREA 0.59 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5175 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.565 1.425 15.7 2.1 ;
      RECT 15.565 2.93 15.62 3.27 ;
      RECT 15.335 1.425 15.565 3.27 ;
      RECT 15.28 1.425 15.335 2.1 ;
      RECT 15.28 2.93 15.335 3.27 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1823 ;
  ANTENNAPARTIALMETALAREA 0.6385 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5387 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.705 1.425 17.005 3.27 ;
      RECT 16.59 1.425 16.705 1.765 ;
      RECT 16.57 2.93 16.705 3.27 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.286 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 1.55 1.84 2.1 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.4107 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3727 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.625 2.48 1.18 3.22 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.265 -0.4 17.16 0.4 ;
      RECT 15.925 -0.4 16.265 1.045 ;
      RECT 14.12 -0.4 15.925 0.4 ;
      RECT 13.78 -0.4 14.12 1.19 ;
      RECT 12.63 -0.4 13.78 0.4 ;
      RECT 12.29 -0.4 12.63 0.575 ;
      RECT 10.54 -0.4 12.29 0.4 ;
      RECT 10.2 -0.4 10.54 0.575 ;
      RECT 8.04 -0.4 10.2 0.4 ;
      RECT 7.7 -0.4 8.04 1.37 ;
      RECT 6.34 -0.4 7.7 0.4 ;
      RECT 6 -0.4 6.34 0.96 ;
      RECT 5.12 -0.4 6 0.44 ;
      RECT 4.695 -0.4 5.12 1.335 ;
      RECT 1.315 -0.4 4.695 0.4 ;
      RECT 0.975 -0.4 1.315 0.575 ;
      RECT 0 -0.4 0.975 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.26 4.64 17.16 5.44 ;
      RECT 15.92 4.08 16.26 5.44 ;
      RECT 14.2 4.64 15.92 5.44 ;
      RECT 13.86 3.68 14.2 5.44 ;
      RECT 11.42 4.64 13.86 5.44 ;
      RECT 11.08 4.08 11.42 5.44 ;
      RECT 8.76 4.64 11.08 5.44 ;
      RECT 7.26 4.08 8.76 5.44 ;
      RECT 4.36 4.64 7.26 5.44 ;
      RECT 4.02 4.465 4.36 5.44 ;
      RECT 1.31 4.64 4.02 5.44 ;
      RECT 0.97 4.465 1.31 5.44 ;
      RECT 0 4.64 0.97 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 16.245 2.095 16.475 2.655 ;
      RECT 16.2 2.425 16.245 2.655 ;
      RECT 15.97 2.425 16.2 3.805 ;
      RECT 14.92 3.575 15.97 3.805 ;
      RECT 14.81 3.575 14.92 4.02 ;
      RECT 14.81 0.85 14.88 1.19 ;
      RECT 14.58 0.85 14.81 4.02 ;
      RECT 14.54 0.85 14.58 1.19 ;
      RECT 14.295 1.59 14.35 2.045 ;
      RECT 14.065 1.59 14.295 3.165 ;
      RECT 14.01 1.59 14.065 2.045 ;
      RECT 13.52 2.935 14.065 3.165 ;
      RECT 13.4 1.815 14.01 2.045 ;
      RECT 13.29 2.935 13.52 3.51 ;
      RECT 13.17 0.91 13.4 2.045 ;
      RECT 12.74 3.28 13.29 3.51 ;
      RECT 13.06 0.91 13.17 1.25 ;
      RECT 12.49 1.815 13.17 2.045 ;
      RECT 12.63 3.28 12.74 3.62 ;
      RECT 12.4 3.28 12.63 4.27 ;
      RECT 12.05 2.46 12.55 2.8 ;
      RECT 12.205 1.63 12.49 2.045 ;
      RECT 12.12 3.93 12.4 4.27 ;
      RECT 12.15 1.63 12.205 1.97 ;
      RECT 11.92 2.46 12.05 3.335 ;
      RECT 11.715 1.685 11.92 3.335 ;
      RECT 11.54 0.635 11.82 0.975 ;
      RECT 11.69 1.27 11.715 3.335 ;
      RECT 11.485 1.27 11.69 1.915 ;
      RECT 11.68 2.68 11.69 3.335 ;
      RECT 10.665 3.105 11.68 3.335 ;
      RECT 11.48 0.635 11.54 1.04 ;
      RECT 9.46 1.27 11.485 1.5 ;
      RECT 11.31 0.69 11.48 1.04 ;
      RECT 11.405 2.205 11.46 2.435 ;
      RECT 11.175 2.205 11.405 2.44 ;
      RECT 9.94 0.81 11.31 1.04 ;
      RECT 10.785 2.21 11.175 2.44 ;
      RECT 10.555 2.04 10.785 2.44 ;
      RECT 10.435 3.105 10.665 3.48 ;
      RECT 9.68 2.04 10.555 2.27 ;
      RECT 10.1 3.25 10.435 3.48 ;
      RECT 9.76 3.25 10.1 3.59 ;
      RECT 9.71 0.63 9.94 1.04 ;
      RECT 9.52 2.6 9.86 2.94 ;
      RECT 8.755 0.63 9.71 0.86 ;
      RECT 9.395 1.735 9.68 2.27 ;
      RECT 9 2.655 9.52 2.885 ;
      RECT 9.23 1.09 9.46 1.5 ;
      RECT 9.34 1.735 9.395 2.075 ;
      RECT 9.06 1.09 9.23 1.43 ;
      RECT 8.77 1.705 9 3.57 ;
      RECT 8.755 1.705 8.77 1.935 ;
      RECT 7.83 3.205 8.77 3.57 ;
      RECT 8.525 0.63 8.755 1.935 ;
      RECT 8.2 2.17 8.54 2.885 ;
      RECT 7.24 1.705 8.525 1.935 ;
      RECT 6.575 2.17 8.2 2.4 ;
      RECT 7.53 2.63 7.87 2.97 ;
      RECT 7.375 2.74 7.53 2.97 ;
      RECT 7.145 2.74 7.375 3.725 ;
      RECT 7.235 1.205 7.24 1.935 ;
      RECT 7.125 1.15 7.235 1.935 ;
      RECT 6.935 3.495 7.145 3.725 ;
      RECT 6.895 0.665 7.125 1.935 ;
      RECT 6.705 3.495 6.935 4.355 ;
      RECT 6.63 0.665 6.895 0.895 ;
      RECT 4.825 4.125 6.705 4.355 ;
      RECT 6.345 1.575 6.575 3.185 ;
      RECT 5.84 1.575 6.345 1.805 ;
      RECT 6.155 2.955 6.345 3.185 ;
      RECT 6.155 3.47 6.21 3.81 ;
      RECT 5.925 2.955 6.155 3.81 ;
      RECT 5.775 2.14 6.115 2.48 ;
      RECT 5.87 3.47 5.925 3.81 ;
      RECT 5.61 1.455 5.84 1.805 ;
      RECT 5.345 2.195 5.775 2.425 ;
      RECT 5.5 1.455 5.61 1.795 ;
      RECT 3.68 1.565 5.5 1.795 ;
      RECT 5.345 3.55 5.4 3.89 ;
      RECT 5.115 2.195 5.345 3.89 ;
      RECT 5.11 2.195 5.115 2.425 ;
      RECT 5.06 3.55 5.115 3.89 ;
      RECT 4.56 2.03 5.11 2.425 ;
      RECT 4.595 3.945 4.825 4.355 ;
      RECT 3.705 3.945 4.595 4.175 ;
      RECT 4.08 0.675 4.42 1.11 ;
      RECT 2.66 0.675 4.08 0.905 ;
      RECT 3.475 2.395 3.705 4.255 ;
      RECT 3.35 1.565 3.68 2.085 ;
      RECT 2.945 2.395 3.475 2.625 ;
      RECT 2.56 4.025 3.475 4.255 ;
      RECT 3.34 1.745 3.35 2.085 ;
      RECT 2.76 3.3 3.1 3.64 ;
      RECT 2.94 1.655 2.945 2.625 ;
      RECT 2.715 1.6 2.94 2.625 ;
      RECT 2.365 3.3 2.76 3.53 ;
      RECT 2.6 1.6 2.715 1.94 ;
      RECT 2.43 0.675 2.66 1.27 ;
      RECT 2.22 3.97 2.56 4.31 ;
      RECT 2.365 0.905 2.43 1.27 ;
      RECT 2.135 0.905 2.365 3.53 ;
      RECT 0.52 4.005 2.22 4.235 ;
      RECT 0.395 1.06 0.52 1.4 ;
      RECT 0.395 3.52 0.52 4.235 ;
      RECT 0.18 1.06 0.395 4.235 ;
      RECT 0.165 1.1 0.18 4.235 ;
  END
END DFFNRX2

MACRO DFFNRX1
  CLASS CORE ;
  FOREIGN DFFNRX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.18 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNRXL ;

  PIN RN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.3139 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3939 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.525 3.34 4.825 3.57 ;
      RECT 4.13 2.95 4.525 3.57 ;
     END
  END RN

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6496 ;
  ANTENNAPARTIALMETALAREA 1.0859 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9131 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.18 2.035 14.41 3.295 ;
      RECT 13.615 2.035 14.18 2.265 ;
      RECT 13.935 3.065 14.18 3.295 ;
      RECT 13.72 3.065 13.935 3.755 ;
      RECT 13.705 3.065 13.72 3.99 ;
      RECT 13.18 3.525 13.705 3.99 ;
      RECT 13.385 1.38 13.615 2.265 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.8885 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6305 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.995 1.355 15 1.85 ;
      RECT 14.735 1.26 14.995 3.98 ;
      RECT 14.66 1.26 14.735 1.85 ;
      RECT 14.44 3.64 14.735 3.98 ;
      RECT 14.59 1.26 14.66 1.75 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.234 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.73 1.78 2.12 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1836 ;
  ANTENNAPARTIALMETALAREA 0.275 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.68 2.67 1.18 3.22 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.33 -0.4 15.18 0.4 ;
      RECT 13.99 -0.4 14.33 0.575 ;
      RECT 12.25 -0.4 13.99 0.4 ;
      RECT 11.91 -0.4 12.25 0.575 ;
      RECT 10.69 -0.4 11.91 0.4 ;
      RECT 10.35 -0.4 10.69 1.31 ;
      RECT 5.975 -0.4 10.35 0.4 ;
      RECT 7.81 1.44 7.92 1.78 ;
      RECT 7.58 1.205 7.81 1.78 ;
      RECT 6.33 1.205 7.58 1.435 ;
      RECT 5.975 1.205 6.33 1.525 ;
      RECT 5.745 -0.4 5.975 1.525 ;
      RECT 4.02 -0.4 5.745 0.4 ;
      RECT 3.68 -0.4 4.02 0.96 ;
      RECT 1.115 -0.4 3.68 0.4 ;
      RECT 0.775 -0.4 1.115 0.575 ;
      RECT 0 -0.4 0.775 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.1 4.64 15.18 5.44 ;
      RECT 13.76 4.465 14.1 5.44 ;
      RECT 12.76 4.64 13.76 5.44 ;
      RECT 12.42 3.62 12.76 5.44 ;
      RECT 10.74 4.64 12.42 5.44 ;
      RECT 10.4 4.07 10.74 5.44 ;
      RECT 8.4 4.64 10.4 5.44 ;
      RECT 7.46 4.07 8.4 5.44 ;
      RECT 4.33 4.64 7.46 5.44 ;
      RECT 3.99 4.465 4.33 5.44 ;
      RECT 1.68 4.64 3.99 5.44 ;
      RECT 1.34 4.465 1.68 5.44 ;
      RECT 0 4.64 1.34 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.42 2.495 13.95 2.835 ;
      RECT 13.145 2.495 13.42 3.14 ;
      RECT 13.08 1.25 13.145 3.14 ;
      RECT 12.845 1.25 13.08 2.795 ;
      RECT 12.79 1.25 12.845 1.55 ;
      RECT 12.45 1.21 12.79 1.55 ;
      RECT 12.455 1.825 12.56 2.11 ;
      RECT 12.225 1.825 12.455 3.295 ;
      RECT 11.925 1.825 12.225 2.055 ;
      RECT 11.48 3.065 12.225 3.295 ;
      RECT 11.695 1.595 11.925 2.055 ;
      RECT 11.39 1.595 11.695 1.825 ;
      RECT 11.14 3.065 11.48 3.94 ;
      RECT 11.39 0.97 11.45 1.31 ;
      RECT 11.11 0.97 11.39 1.825 ;
      RECT 11.325 2.14 11.38 2.48 ;
      RECT 11.04 2.14 11.325 2.505 ;
      RECT 10.54 1.595 11.11 1.825 ;
      RECT 9.915 2.275 11.04 2.505 ;
      RECT 10.255 1.595 10.54 2.045 ;
      RECT 10.2 1.705 10.255 2.045 ;
      RECT 9.915 4 10.03 4.34 ;
      RECT 9.905 2.275 9.915 4.34 ;
      RECT 9.685 2.02 9.905 4.34 ;
      RECT 9.675 2.02 9.685 4.285 ;
      RECT 9.225 2.02 9.675 2.25 ;
      RECT 9.22 0.65 9.56 0.99 ;
      RECT 9.225 1.23 9.28 1.57 ;
      RECT 8.605 2.5 9.26 2.84 ;
      RECT 8.995 1.23 9.225 2.25 ;
      RECT 8.605 0.675 9.22 0.905 ;
      RECT 8.94 1.23 8.995 1.57 ;
      RECT 8.375 0.675 8.605 3.33 ;
      RECT 6.545 0.675 8.375 0.905 ;
      RECT 8.12 3.1 8.375 3.33 ;
      RECT 7.78 3.1 8.12 3.44 ;
      RECT 8.005 2.02 8.06 2.41 ;
      RECT 7.72 2.02 8.005 2.415 ;
      RECT 6.645 2.18 7.72 2.415 ;
      RECT 7.295 2.705 7.525 3.825 ;
      RECT 7.165 3.595 7.295 3.825 ;
      RECT 6.935 3.595 7.165 4.365 ;
      RECT 4.79 4.135 6.935 4.365 ;
      RECT 6.415 1.825 6.645 3.385 ;
      RECT 6.205 0.635 6.545 0.975 ;
      RECT 5.38 1.825 6.415 2.055 ;
      RECT 6.11 3.155 6.415 3.385 ;
      RECT 5.88 3.155 6.11 3.82 ;
      RECT 5.76 2.44 6.1 2.78 ;
      RECT 5.77 3.48 5.88 3.82 ;
      RECT 5.355 2.495 5.76 2.725 ;
      RECT 5.355 3.48 5.41 3.82 ;
      RECT 5.37 1.655 5.38 2.055 ;
      RECT 5.15 1.18 5.37 2.055 ;
      RECT 5.125 2.435 5.355 3.82 ;
      RECT 5.14 1.18 5.15 1.885 ;
      RECT 3.57 1.655 5.14 1.885 ;
      RECT 4.92 2.435 5.125 2.665 ;
      RECT 5.07 3.48 5.125 3.82 ;
      RECT 4.555 2.12 4.92 2.665 ;
      RECT 4.565 0.77 4.87 1.11 ;
      RECT 4.56 3.945 4.79 4.365 ;
      RECT 4.335 0.77 4.565 1.42 ;
      RECT 3.675 3.945 4.56 4.175 ;
      RECT 2.53 1.19 4.335 1.42 ;
      RECT 3.465 2.935 3.675 4.355 ;
      RECT 3.23 1.655 3.57 2.08 ;
      RECT 3.445 2.395 3.465 4.355 ;
      RECT 3.235 2.395 3.445 3.165 ;
      RECT 2.145 4.125 3.445 4.355 ;
      RECT 2.905 2.395 3.235 2.625 ;
      RECT 2.775 3.48 3.11 3.84 ;
      RECT 2.845 2.105 2.905 2.625 ;
      RECT 2.675 1.94 2.845 2.625 ;
      RECT 2.545 2.855 2.775 3.84 ;
      RECT 2.615 1.94 2.675 2.335 ;
      RECT 2.38 2.855 2.545 3.085 ;
      RECT 2.38 1.16 2.53 1.5 ;
      RECT 2.19 1.16 2.38 3.085 ;
      RECT 2.15 1.22 2.19 3.085 ;
      RECT 1.915 3.745 2.145 4.355 ;
      RECT 0.845 3.745 1.915 3.975 ;
      RECT 0.505 3.52 0.845 3.975 ;
      RECT 0.39 1.15 0.52 1.49 ;
      RECT 0.39 3.52 0.505 3.75 ;
      RECT 0.18 1.15 0.39 3.75 ;
      RECT 0.16 1.26 0.18 3.75 ;
  END
END DFFNRX1

MACRO DFFNXL
  CLASS CORE ;
  FOREIGN DFFNXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.22 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6624 ;
  ANTENNAPARTIALMETALAREA 0.9146 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2118 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.7 1.2 11.04 3.79 ;
      RECT 10.6 3.45 10.7 3.79 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.4564 ;
  ANTENNAPARTIALMETALAREA 1.1582 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.2947 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.115 0.865 10.345 3.42 ;
      RECT 10.04 0.865 10.115 1.285 ;
      RECT 9.29 3.19 10.115 3.42 ;
      RECT 9.83 0.865 10.04 1.095 ;
      RECT 9.3 0.745 9.83 1.095 ;
      RECT 8.95 3.19 9.29 3.53 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.345 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.305 1.675 1.84 2.32 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3156 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1925 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.645 2.63 1.18 3.22 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.46 -0.4 11.22 0.4 ;
      RECT 10.12 -0.4 10.46 0.575 ;
      RECT 8.88 -0.4 10.12 0.4 ;
      RECT 8.54 -0.4 8.88 0.575 ;
      RECT 6.4 -0.4 8.54 0.4 ;
      RECT 6.06 -0.4 6.4 1.555 ;
      RECT 4.07 -0.4 6.06 0.4 ;
      RECT 3.73 -0.4 4.07 1.15 ;
      RECT 1.265 -0.4 3.73 0.4 ;
      RECT 0.925 -0.4 1.265 0.575 ;
      RECT 0 -0.4 0.925 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.18 4.64 11.22 5.44 ;
      RECT 9.84 4.41 10.18 5.44 ;
      RECT 8.47 4.64 9.84 5.44 ;
      RECT 8.13 4.465 8.47 5.44 ;
      RECT 5.795 4.64 8.13 5.44 ;
      RECT 5.455 4.465 5.795 5.44 ;
      RECT 1.485 4.64 5.455 5.44 ;
      RECT 1.145 4.41 1.485 5.44 ;
      RECT 0 4.64 1.145 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.805 2.005 9.87 2.375 ;
      RECT 9.68 1.47 9.805 2.945 ;
      RECT 9.575 1.46 9.68 2.945 ;
      RECT 9.34 1.46 9.575 1.8 ;
      RECT 8.4 2.715 9.575 2.945 ;
      RECT 8.915 2.105 9.255 2.445 ;
      RECT 9.175 4.06 9.23 4.4 ;
      RECT 8.89 3.97 9.175 4.4 ;
      RECT 8.88 2.105 8.915 2.335 ;
      RECT 8.4 3.97 8.89 4.2 ;
      RECT 8.65 1.44 8.88 2.335 ;
      RECT 7.55 1.44 8.65 1.835 ;
      RECT 8.35 2.715 8.4 4.2 ;
      RECT 8.17 2.18 8.35 4.2 ;
      RECT 8.01 2.18 8.17 2.945 ;
      RECT 7.76 0.835 8.1 1.175 ;
      RECT 6.94 0.945 7.76 1.175 ;
      RECT 7.32 1.44 7.55 4.15 ;
      RECT 7.26 3.92 7.32 4.15 ;
      RECT 6.92 3.92 7.26 4.26 ;
      RECT 6.98 1.84 7.09 3.16 ;
      RECT 6.94 1.84 6.98 3.615 ;
      RECT 6.75 0.945 6.94 3.615 ;
      RECT 6.71 0.945 6.75 2.07 ;
      RECT 6.27 3.385 6.75 3.615 ;
      RECT 5.6 1.84 6.71 2.07 ;
      RECT 6.31 2.38 6.42 2.72 ;
      RECT 6.08 2.38 6.31 3.135 ;
      RECT 6.04 3.385 6.27 4.235 ;
      RECT 5.8 2.905 6.08 3.135 ;
      RECT 3.59 4.005 6.04 4.235 ;
      RECT 5.57 2.905 5.8 3.775 ;
      RECT 5.33 1.21 5.6 2.07 ;
      RECT 4.76 3.545 5.57 3.775 ;
      RECT 5.26 1.21 5.33 3.12 ;
      RECT 5.1 1.84 5.26 3.12 ;
      RECT 4.99 2.78 5.1 3.12 ;
      RECT 4.815 0.83 4.87 1.17 ;
      RECT 4.76 0.83 4.815 2.47 ;
      RECT 4.585 0.83 4.76 3.775 ;
      RECT 4.53 0.83 4.585 1.17 ;
      RECT 4.49 2.22 4.585 3.775 ;
      RECT 3.58 2.22 4.49 2.56 ;
      RECT 4.015 1.485 4.355 1.825 ;
      RECT 3.375 1.595 4.015 1.825 ;
      RECT 3.48 3.95 3.59 4.29 ;
      RECT 3.25 3.72 3.48 4.29 ;
      RECT 3.295 1.195 3.375 1.825 ;
      RECT 3.295 3.15 3.35 3.49 ;
      RECT 3.065 1.195 3.295 3.49 ;
      RECT 2.49 3.72 3.25 3.95 ;
      RECT 2.71 1.195 3.065 1.48 ;
      RECT 3.01 3.15 3.065 3.49 ;
      RECT 2.03 4.18 2.895 4.41 ;
      RECT 2.37 1.14 2.71 1.48 ;
      RECT 2.43 1.845 2.49 3.95 ;
      RECT 2.26 1.735 2.43 3.95 ;
      RECT 2.09 1.735 2.26 2.075 ;
      RECT 1.8 3.605 2.03 4.41 ;
      RECT 0.65 3.605 1.8 3.835 ;
      RECT 0.415 3.455 0.65 3.835 ;
      RECT 0.415 1.2 0.53 1.54 ;
      RECT 0.19 1.2 0.415 3.835 ;
      RECT 0.185 1.255 0.19 3.835 ;
  END
END DFFNXL

MACRO DFFNX4
  CLASS CORE ;
  FOREIGN DFFNX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2684 ;
  ANTENNAPARTIALMETALAREA 0.7481 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5705 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.01 1.82 15.04 3.22 ;
      RECT 14.965 1.29 15.01 3.22 ;
      RECT 14.945 1.29 14.965 3.225 ;
      RECT 14.67 1.29 14.945 3.28 ;
      RECT 14.66 1.82 14.67 3.28 ;
      RECT 14.605 2.94 14.66 3.28 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2684 ;
  ANTENNAPARTIALMETALAREA 0.7371 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5387 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.72 1.29 13.73 1.85 ;
      RECT 13.675 1.29 13.72 3.22 ;
      RECT 13.665 1.29 13.675 3.225 ;
      RECT 13.39 1.29 13.665 3.28 ;
      RECT 13.34 1.82 13.39 3.28 ;
      RECT 13.325 2.94 13.34 3.28 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.234 ;
  ANTENNAPARTIALMETALAREA 0.3111 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.6059 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.365 2.4 1.595 3.185 ;
      RECT 1.125 2.89 1.365 3.185 ;
      RECT 1.105 2.955 1.125 3.185 ;
      RECT 0.875 2.955 1.105 3.195 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.4788 ;
  ANTENNAPARTIALMETALAREA 0.2863 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5635 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.925 1.845 1.765 2.075 ;
      RECT 0.695 1.845 0.925 2.25 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.65 -0.4 15.84 0.4 ;
      RECT 15.31 -0.4 15.65 0.965 ;
      RECT 14.37 -0.4 15.31 0.4 ;
      RECT 14.03 -0.4 14.37 0.965 ;
      RECT 13.09 -0.4 14.03 0.4 ;
      RECT 12.75 -0.4 13.09 0.965 ;
      RECT 11.61 -0.4 12.75 0.4 ;
      RECT 11.27 -0.4 11.61 0.575 ;
      RECT 8.91 -0.4 11.27 0.4 ;
      RECT 8.57 -0.4 8.91 1.28 ;
      RECT 6.35 -0.4 8.57 0.4 ;
      RECT 6.01 -0.4 6.35 1.435 ;
      RECT 3.925 -0.4 6.01 0.4 ;
      RECT 3.585 -0.4 3.925 1.375 ;
      RECT 1.32 -0.4 3.585 0.4 ;
      RECT 0.98 -0.4 1.32 0.575 ;
      RECT 0 -0.4 0.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.585 4.64 15.84 5.44 ;
      RECT 15.245 4.075 15.585 5.44 ;
      RECT 14.305 4.64 15.245 5.44 ;
      RECT 13.965 4.075 14.305 5.44 ;
      RECT 13.025 4.64 13.965 5.44 ;
      RECT 12.685 4.075 13.025 5.44 ;
      RECT 11.46 4.64 12.685 5.44 ;
      RECT 11.09 4.4 11.46 5.44 ;
      RECT 8.88 4.64 11.09 5.44 ;
      RECT 8.54 4.09 8.88 5.44 ;
      RECT 6.265 4.64 8.54 5.44 ;
      RECT 5.925 4.465 6.265 5.44 ;
      RECT 4 4.64 5.925 5.44 ;
      RECT 3.66 4.465 4 5.44 ;
      RECT 1.4 4.64 3.66 5.44 ;
      RECT 1.06 4.465 1.4 5.44 ;
      RECT 0 4.64 1.06 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.325 2.29 15.555 3.755 ;
      RECT 12.995 3.525 15.325 3.755 ;
      RECT 12.765 1.265 12.995 3.755 ;
      RECT 12.37 1.265 12.765 1.495 ;
      RECT 12.24 3.42 12.765 3.755 ;
      RECT 12.285 2.29 12.515 3.045 ;
      RECT 12.03 1.13 12.37 1.495 ;
      RECT 10.97 2.815 12.285 3.045 ;
      RECT 11.9 3.42 12.24 3.76 ;
      RECT 11.43 1.265 12.03 1.495 ;
      RECT 11.2 1.265 11.43 2.58 ;
      RECT 10.74 0.995 10.97 3.855 ;
      RECT 9.625 0.995 10.74 1.225 ;
      RECT 10.16 3.625 10.74 3.855 ;
      RECT 10.275 1.495 10.505 2.905 ;
      RECT 9.92 2.675 10.275 2.905 ;
      RECT 9.82 3.625 10.16 3.99 ;
      RECT 9.81 2.595 9.92 2.935 ;
      RECT 7.6 3.625 9.82 3.855 ;
      RECT 9.58 2.595 9.81 3.335 ;
      RECT 9.395 0.995 9.625 1.825 ;
      RECT 7.59 3.105 9.58 3.335 ;
      RECT 7.685 1.595 9.395 1.825 ;
      RECT 8.82 2.14 9.11 2.48 ;
      RECT 8.3 2.065 8.82 2.48 ;
      RECT 6.615 2.065 8.3 2.295 ;
      RECT 7.63 1.33 7.685 1.825 ;
      RECT 7.455 1.275 7.63 1.825 ;
      RECT 7.315 3.625 7.6 4.08 ;
      RECT 7.25 2.53 7.59 3.335 ;
      RECT 7.29 1.275 7.455 1.615 ;
      RECT 7.26 3.74 7.315 4.08 ;
      RECT 5.48 3.105 7.25 3.335 ;
      RECT 6.205 1.67 6.615 2.36 ;
      RECT 5.78 1.67 6.205 1.9 ;
      RECT 5.55 0.935 5.78 1.9 ;
      RECT 4.685 0.935 5.55 1.165 ;
      RECT 5.425 3.06 5.48 3.4 ;
      RECT 5.32 3.06 5.425 4.175 ;
      RECT 5.195 1.42 5.32 4.175 ;
      RECT 5.09 1.42 5.195 3.425 ;
      RECT 3.205 3.945 5.195 4.175 ;
      RECT 4.685 2.72 4.705 3.71 ;
      RECT 4.475 0.935 4.685 3.71 ;
      RECT 4.455 0.935 4.475 2.95 ;
      RECT 4.31 1.13 4.455 1.47 ;
      RECT 3.365 2.61 4.455 2.95 ;
      RECT 3.8 1.89 4.14 2.23 ;
      RECT 3.095 1.945 3.8 2.175 ;
      RECT 2.975 3.945 3.205 4.235 ;
      RECT 3.065 1.375 3.095 2.175 ;
      RECT 2.835 1.375 3.065 3.515 ;
      RECT 2.165 4.005 2.975 4.235 ;
      RECT 1.78 0.675 2.97 0.905 ;
      RECT 2.54 1.375 2.835 1.605 ;
      RECT 2.665 3.285 2.835 3.515 ;
      RECT 2.435 3.285 2.665 3.65 ;
      RECT 2.255 1.24 2.54 1.605 ;
      RECT 2.165 1.92 2.305 2.995 ;
      RECT 2.2 1.24 2.255 1.58 ;
      RECT 2.075 1.92 2.165 4.235 ;
      RECT 1.935 2.765 2.075 4.235 ;
      RECT 1.55 0.675 1.78 1.395 ;
      RECT 0.56 1.165 1.55 1.395 ;
      RECT 0.43 1.165 0.56 1.53 ;
      RECT 0.43 2.9 0.54 4.18 ;
      RECT 0.275 1.165 0.43 4.18 ;
      RECT 0.22 1.19 0.275 4.18 ;
      RECT 0.2 1.245 0.22 4.18 ;
  END
END DFFNX4

MACRO DFFNX2
  CLASS CORE ;
  FOREIGN DFFNX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.81 ;
  ANTENNAPARTIALMETALAREA 0.6532 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0581 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.755 1.355 12.985 3.33 ;
      RECT 12.68 1.355 12.755 1.845 ;
      RECT 12.7 3.1 12.755 3.33 ;
      RECT 12.36 3.1 12.7 3.44 ;
      RECT 12.58 1.355 12.68 1.695 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8456 ;
  ANTENNAPARTIALMETALAREA 0.9031 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9644 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.505 0.7 11.56 1.04 ;
      RECT 11.22 0.7 11.505 1.08 ;
      RECT 10.865 0.85 11.22 1.08 ;
      RECT 11.08 2.88 11.16 3.22 ;
      RECT 10.865 2.635 11.08 3.22 ;
      RECT 10.7 0.85 10.865 3.22 ;
      RECT 10.635 0.85 10.7 3.165 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.162 ;
  ANTENNAPARTIALMETALAREA 0.3507 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4151 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.405 1.825 2.24 ;
      RECT 1.325 1.405 1.46 1.745 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.228 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.06 1.18 2.66 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.48 -0.4 13.86 0.4 ;
      RECT 13.14 -0.4 13.48 0.575 ;
      RECT 12.36 -0.4 13.14 0.4 ;
      RECT 12.02 -0.4 12.36 0.575 ;
      RECT 10.76 -0.4 12.02 0.4 ;
      RECT 10.42 -0.4 10.76 0.575 ;
      RECT 8.8 -0.4 10.42 0.4 ;
      RECT 8.46 -0.4 8.8 1.27 ;
      RECT 6.185 -0.4 8.46 0.4 ;
      RECT 5.845 -0.4 6.185 1.44 ;
      RECT 4.02 -0.4 5.845 0.4 ;
      RECT 3.68 -0.4 4.02 1.285 ;
      RECT 1.285 -0.4 3.68 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.26 4.64 13.86 5.44 ;
      RECT 12.92 4.465 13.26 5.44 ;
      RECT 11.92 4.64 12.92 5.44 ;
      RECT 11.58 4.465 11.92 5.44 ;
      RECT 9.94 4.64 11.58 5.44 ;
      RECT 8.19 4.465 9.94 5.44 ;
      RECT 5.87 4.64 8.19 5.44 ;
      RECT 5.53 4.465 5.87 5.44 ;
      RECT 4.53 4.64 5.53 5.44 ;
      RECT 4.19 4.465 4.53 5.44 ;
      RECT 1.34 4.64 4.19 5.44 ;
      RECT 1 4.41 1.34 5.44 ;
      RECT 0 4.64 1 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.435 4.02 12.49 4.36 ;
      RECT 12.15 3.995 12.435 4.36 ;
      RECT 12.125 3.995 12.15 4.225 ;
      RECT 11.895 1.535 12.125 4.225 ;
      RECT 11.22 1.535 11.895 1.765 ;
      RECT 11.16 3.995 11.895 4.225 ;
      RECT 11.435 2.275 11.665 3.68 ;
      RECT 9.975 3.45 11.435 3.68 ;
      RECT 11.05 3.995 11.16 4.37 ;
      RECT 10.82 3.91 11.05 4.37 ;
      RECT 9.64 3.91 10.82 4.14 ;
      RECT 9.745 1.775 9.975 3.68 ;
      RECT 9.6 1.775 9.745 2.005 ;
      RECT 9.03 3.415 9.745 3.68 ;
      RECT 9.37 1.145 9.6 2.005 ;
      RECT 9.11 2.35 9.45 2.69 ;
      RECT 9.26 1.145 9.37 1.795 ;
      RECT 8.13 1.565 9.26 1.795 ;
      RECT 8.195 2.405 9.11 2.635 ;
      RECT 8.92 3.36 9.03 3.7 ;
      RECT 8.69 3.36 8.92 3.96 ;
      RECT 7.155 3.73 8.69 3.96 ;
      RECT 7.965 2.405 8.195 3.13 ;
      RECT 7.9 1.16 8.13 1.795 ;
      RECT 7.3 2.9 7.965 3.13 ;
      RECT 7.52 1.16 7.9 1.39 ;
      RECT 7.18 1.05 7.52 1.39 ;
      RECT 7.21 2.82 7.3 3.16 ;
      RECT 6.98 1.77 7.21 3.16 ;
      RECT 6.925 3.44 7.155 4.275 ;
      RECT 5.39 1.77 6.98 2 ;
      RECT 6.96 2.82 6.98 3.16 ;
      RECT 6.33 2.93 6.96 3.16 ;
      RECT 5.86 2.245 6.61 2.475 ;
      RECT 6.1 2.93 6.33 4.235 ;
      RECT 3.595 4.005 6.1 4.235 ;
      RECT 5.63 2.245 5.86 3.755 ;
      RECT 4.695 3.525 5.63 3.755 ;
      RECT 5.39 1.095 5.445 1.435 ;
      RECT 5.38 1.095 5.39 2 ;
      RECT 5.33 1.095 5.38 2.91 ;
      RECT 5.15 1.095 5.33 2.965 ;
      RECT 5.105 1.095 5.15 1.435 ;
      RECT 4.99 2.625 5.15 2.965 ;
      RECT 4.685 2.27 4.695 3.755 ;
      RECT 4.465 0.965 4.685 3.755 ;
      RECT 4.455 0.965 4.465 2.58 ;
      RECT 3.925 2.17 4.455 2.5 ;
      RECT 3.355 1.555 4.18 1.785 ;
      RECT 3.585 2.17 3.925 2.51 ;
      RECT 3.365 3.695 3.595 4.235 ;
      RECT 2.895 3.695 3.365 3.925 ;
      RECT 3.125 1.545 3.355 3.43 ;
      RECT 2.97 1.545 3.125 1.785 ;
      RECT 2.74 0.92 2.97 1.785 ;
      RECT 2.665 2.82 2.895 3.925 ;
      RECT 1.98 4.18 2.84 4.41 ;
      RECT 2.66 0.92 2.74 1.15 ;
      RECT 2.375 2.82 2.665 3.05 ;
      RECT 2.32 0.81 2.66 1.15 ;
      RECT 2.375 1.38 2.43 1.72 ;
      RECT 2.145 1.38 2.375 3.05 ;
      RECT 2.09 1.38 2.145 1.72 ;
      RECT 1.75 3.605 1.98 4.41 ;
      RECT 0.79 3.605 1.75 3.835 ;
      RECT 0.57 3.02 0.79 3.835 ;
      RECT 0.39 1.34 0.57 3.835 ;
      RECT 0.34 1.34 0.39 3.31 ;
      RECT 0.18 1.34 0.34 1.68 ;
  END
END DFFNX2

MACRO DFFNX1
  CLASS CORE ;
  FOREIGN DFFNX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.22 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFNXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.936 ;
  ANTENNAPARTIALMETALAREA 0.9486 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3178 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.7 1.19 11.04 3.88 ;
      RECT 10.6 3.54 10.7 3.88 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5214 ;
  ANTENNAPARTIALMETALAREA 1.1537 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.115 0.865 10.345 3.42 ;
      RECT 9.64 0.865 10.115 1.095 ;
      RECT 9.23 3.19 10.115 3.42 ;
      RECT 9.3 0.69 9.64 1.095 ;
      RECT 8.89 3.19 9.23 3.53 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1314 ;
  ANTENNAPARTIALMETALAREA 0.3245 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.29 1.82 1.84 2.41 ;
     END
  END D

  PIN CKN
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.2862 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.645 2.685 1.18 3.22 ;
     END
  END CKN

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.46 -0.4 11.22 0.4 ;
      RECT 10.12 -0.4 10.46 0.575 ;
      RECT 8.88 -0.4 10.12 0.4 ;
      RECT 8.54 -0.4 8.88 0.575 ;
      RECT 6.44 -0.4 8.54 0.4 ;
      RECT 6.1 -0.4 6.44 1.46 ;
      RECT 4.07 -0.4 6.1 0.4 ;
      RECT 3.73 -0.4 4.07 1.15 ;
      RECT 1.305 -0.4 3.73 0.4 ;
      RECT 0.965 -0.4 1.305 0.575 ;
      RECT 0 -0.4 0.965 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.18 4.64 11.22 5.44 ;
      RECT 9.84 4.41 10.18 5.44 ;
      RECT 8.47 4.64 9.84 5.44 ;
      RECT 8.13 4.465 8.47 5.44 ;
      RECT 5.8 4.64 8.13 5.44 ;
      RECT 4.52 4.465 5.8 5.44 ;
      RECT 1.035 4.64 4.52 5.44 ;
      RECT 0.695 4.41 1.035 5.44 ;
      RECT 0 4.64 0.695 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.64 1.47 9.87 2.76 ;
      RECT 9.34 1.47 9.64 1.81 ;
      RECT 8.4 2.53 9.64 2.76 ;
      RECT 8.88 2.065 9.255 2.295 ;
      RECT 8.89 3.99 9.23 4.37 ;
      RECT 8.4 3.99 8.89 4.22 ;
      RECT 8.65 1.44 8.88 2.295 ;
      RECT 7.55 1.44 8.65 1.835 ;
      RECT 8.35 2.53 8.4 4.22 ;
      RECT 8.17 2.18 8.35 4.22 ;
      RECT 8.065 2.18 8.17 2.76 ;
      RECT 6.94 0.67 8.1 0.9 ;
      RECT 8.01 2.18 8.065 2.52 ;
      RECT 7.32 1.44 7.55 4.23 ;
      RECT 7.21 4 7.32 4.23 ;
      RECT 6.87 4 7.21 4.34 ;
      RECT 6.865 2.82 7.09 3.16 ;
      RECT 6.865 0.67 6.94 1.995 ;
      RECT 6.71 0.67 6.865 3.615 ;
      RECT 6.635 1.765 6.71 3.615 ;
      RECT 5.555 1.84 6.635 2.07 ;
      RECT 6.27 3.385 6.635 3.615 ;
      RECT 6.135 2.38 6.365 3.135 ;
      RECT 6.04 3.385 6.27 4.235 ;
      RECT 5.8 2.905 6.135 3.135 ;
      RECT 3.59 4.005 6.04 4.235 ;
      RECT 5.57 2.905 5.8 3.775 ;
      RECT 5.555 1.17 5.61 1.51 ;
      RECT 4.76 3.545 5.57 3.775 ;
      RECT 5.315 1.17 5.555 2.07 ;
      RECT 5.315 2.79 5.33 3.13 ;
      RECT 5.27 1.17 5.315 3.13 ;
      RECT 5.085 1.84 5.27 3.13 ;
      RECT 4.99 2.79 5.085 3.13 ;
      RECT 4.815 0.83 4.87 1.17 ;
      RECT 4.76 0.83 4.815 2.47 ;
      RECT 4.585 0.83 4.76 3.775 ;
      RECT 4.53 0.83 4.585 1.17 ;
      RECT 4.49 2.2 4.585 3.775 ;
      RECT 3.58 2.2 4.49 2.54 ;
      RECT 4.015 1.425 4.355 1.765 ;
      RECT 3.295 1.425 4.015 1.655 ;
      RECT 3.485 3.95 3.59 4.29 ;
      RECT 3.25 3.72 3.485 4.29 ;
      RECT 3.295 3.15 3.35 3.49 ;
      RECT 3.065 1.17 3.295 3.49 ;
      RECT 2.375 3.72 3.25 3.95 ;
      RECT 2.71 1.17 3.065 1.4 ;
      RECT 3.01 3.15 3.065 3.49 ;
      RECT 1.765 4.18 2.895 4.41 ;
      RECT 2.37 1.06 2.71 1.4 ;
      RECT 2.145 1.685 2.375 3.95 ;
      RECT 1.535 3.605 1.765 4.41 ;
      RECT 0.65 3.605 1.535 3.835 ;
      RECT 0.415 3.455 0.65 3.835 ;
      RECT 0.415 1.095 0.53 1.435 ;
      RECT 0.19 1.095 0.415 3.835 ;
      RECT 0.185 1.15 0.19 3.835 ;
  END
END DFFNX1

MACRO DFFHQXL
  CLASS CORE ;
  FOREIGN DFFHQXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 1.2275 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.3159 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.345 0.74 10.435 3.53 ;
      RECT 10.205 0.74 10.345 3.755 ;
      RECT 9.59 0.74 10.205 0.97 ;
      RECT 10.115 3.19 10.205 3.755 ;
      RECT 9.05 3.19 10.115 3.53 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.3483 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3144 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.41 1.82 1.84 2.63 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2484 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.745 2.08 1.105 2.77 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.17 -0.4 10.56 0.4 ;
      RECT 8.83 -0.4 9.17 0.575 ;
      RECT 6.315 -0.4 8.83 0.4 ;
      RECT 6.085 -0.4 6.315 1.46 ;
      RECT 4.015 -0.4 6.085 0.4 ;
      RECT 3.785 -0.4 4.015 1.15 ;
      RECT 1.35 -0.4 3.785 0.4 ;
      RECT 1.01 -0.4 1.35 0.575 ;
      RECT 0 -0.4 1.01 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.63 4.64 10.56 5.44 ;
      RECT 8.29 4.465 8.63 5.44 ;
      RECT 5.795 4.64 8.29 5.44 ;
      RECT 5.455 4.465 5.795 5.44 ;
      RECT 1.815 4.64 5.455 5.44 ;
      RECT 1.475 4.465 1.815 5.44 ;
      RECT 0 4.64 1.475 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.925 1.46 9.97 1.8 ;
      RECT 9.695 1.46 9.925 2.96 ;
      RECT 9.63 1.46 9.695 1.8 ;
      RECT 8.64 2.73 9.695 2.96 ;
      RECT 9.235 2.04 9.465 2.38 ;
      RECT 9.09 4.115 9.39 4.345 ;
      RECT 9.17 2.04 9.235 2.27 ;
      RECT 8.94 1.605 9.17 2.27 ;
      RECT 8.86 4.005 9.09 4.345 ;
      RECT 7.955 1.605 8.94 1.835 ;
      RECT 8.64 4.005 8.86 4.235 ;
      RECT 8.41 2.18 8.64 4.235 ;
      RECT 8.3 2.18 8.41 2.52 ;
      RECT 6.775 0.875 8.39 1.105 ;
      RECT 7.725 1.37 7.955 4.375 ;
      RECT 7.03 4.145 7.725 4.375 ;
      RECT 7.265 1.715 7.495 3.915 ;
      RECT 7.235 1.715 7.265 1.945 ;
      RECT 6.595 3.685 7.265 3.915 ;
      RECT 7.005 1.345 7.235 1.945 ;
      RECT 6.805 2.225 7.035 3.455 ;
      RECT 6.775 2.225 6.805 2.455 ;
      RECT 6.135 3.225 6.805 3.455 ;
      RECT 6.545 0.875 6.775 2.455 ;
      RECT 6.365 3.685 6.595 4.14 ;
      RECT 5.56 1.765 6.545 1.995 ;
      RECT 5.675 2.745 6.42 2.975 ;
      RECT 5.905 3.225 6.135 4.235 ;
      RECT 2.375 4.005 5.905 4.235 ;
      RECT 5.445 2.745 5.675 3.775 ;
      RECT 5.365 1.17 5.57 1.51 ;
      RECT 4.68 3.545 5.445 3.775 ;
      RECT 5.275 0.63 5.365 1.51 ;
      RECT 5.215 0.63 5.275 1.94 ;
      RECT 5.135 0.63 5.215 3.13 ;
      RECT 5.045 1.225 5.135 3.13 ;
      RECT 4.985 1.71 5.045 3.13 ;
      RECT 4.68 0.81 4.815 1.465 ;
      RECT 4.585 0.81 4.68 3.775 ;
      RECT 4.45 1.235 4.585 3.775 ;
      RECT 4.395 2.185 4.45 3.775 ;
      RECT 3.92 2.185 4.395 2.415 ;
      RECT 3.295 1.515 4.22 1.745 ;
      RECT 3.58 2.13 3.92 2.47 ;
      RECT 3.065 0.805 3.295 3.68 ;
      RECT 2.37 0.805 3.065 1.035 ;
      RECT 2.145 1.41 2.375 4.235 ;
      RECT 1.055 3.135 2.145 3.365 ;
      RECT 0.715 3.025 1.055 3.365 ;
      RECT 0.415 1.41 0.75 1.75 ;
      RECT 0.415 3.025 0.715 3.255 ;
      RECT 0.185 1.41 0.415 3.255 ;
  END
END DFFHQXL

MACRO DFFHQX4
  CLASS CORE ;
  FOREIGN DFFHQX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.52 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFHQXL ;

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.6038 ;
  ANTENNAPARTIALMETALAREA 1.0608 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6252 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.62 1.82 13.72 3.22 ;
      RECT 13.54 0.835 13.62 3.22 ;
      RECT 13.34 0.835 13.54 3.675 ;
      RECT 13.28 0.835 13.34 1.645 ;
      RECT 13.2 2.865 13.34 3.675 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.234 ;
  ANTENNAPARTIALMETALAREA 0.2869 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.415 2.605 1.84 3.28 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.414 ;
  ANTENNAPARTIALMETALAREA 0.2109 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9752 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.62 2.2 1.105 2.635 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.34 -0.4 14.52 0.4 ;
      RECT 14 -0.4 14.34 1.015 ;
      RECT 12.86 -0.4 14 0.4 ;
      RECT 12.52 -0.4 12.86 0.575 ;
      RECT 11.56 -0.4 12.52 0.4 ;
      RECT 11.22 -0.4 11.56 1.25 ;
      RECT 9.345 -0.4 11.22 0.4 ;
      RECT 9.115 -0.4 9.345 1.27 ;
      RECT 6.205 -0.4 9.115 0.4 ;
      RECT 5.975 -0.4 6.205 1.37 ;
      RECT 3.82 -0.4 5.975 0.4 ;
      RECT 3.48 -0.4 3.82 1.27 ;
      RECT 1.3 -0.4 3.48 0.4 ;
      RECT 0.96 -0.4 1.3 0.575 ;
      RECT 0 -0.4 0.96 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.3 4.64 14.52 5.44 ;
      RECT 13.96 4.465 14.3 5.44 ;
      RECT 12.78 4.64 13.96 5.44 ;
      RECT 12.44 4.465 12.78 5.44 ;
      RECT 11.4 4.64 12.44 5.44 ;
      RECT 9.65 4.465 11.4 5.44 ;
      RECT 6.13 4.64 9.65 5.44 ;
      RECT 5.79 4.465 6.13 5.44 ;
      RECT 4.065 4.64 5.79 5.44 ;
      RECT 3.725 4.465 4.065 5.44 ;
      RECT 1.37 4.64 3.725 5.44 ;
      RECT 1.03 4.465 1.37 5.44 ;
      RECT 0 4.64 1.03 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.305 2.065 12.31 3.81 ;
      RECT 12.08 1.195 12.305 3.81 ;
      RECT 12.075 1.195 12.08 2.43 ;
      RECT 11.82 3.47 12.08 3.81 ;
      RECT 11.385 2.2 12.075 2.43 ;
      RECT 11.155 2.87 11.84 3.1 ;
      RECT 10.925 1.5 11.155 3.965 ;
      RECT 10.2 1.5 10.925 1.73 ;
      RECT 10.125 3.735 10.925 3.965 ;
      RECT 10.465 1.96 10.695 3.235 ;
      RECT 8.42 1.96 10.465 2.19 ;
      RECT 9.66 3.005 10.465 3.235 ;
      RECT 10.005 2.425 10.235 2.77 ;
      RECT 9.86 0.965 10.2 1.73 ;
      RECT 9.895 3.735 10.125 4.03 ;
      RECT 9.2 2.54 10.005 2.77 ;
      RECT 7.83 3.8 9.895 4.03 ;
      RECT 9.855 1.075 9.86 1.73 ;
      RECT 8.885 1.5 9.855 1.73 ;
      RECT 9.43 3.005 9.66 3.57 ;
      RECT 6.77 3.34 9.43 3.57 ;
      RECT 8.97 2.54 9.2 3.11 ;
      RECT 7.5 2.88 8.97 3.11 ;
      RECT 8.655 1.05 8.885 1.73 ;
      RECT 7.96 2.42 8.74 2.65 ;
      RECT 7.36 1.05 8.655 1.28 ;
      RECT 8.19 1.515 8.42 2.19 ;
      RECT 7.125 1.515 8.19 1.745 ;
      RECT 7.73 2.035 7.96 2.65 ;
      RECT 7.49 3.8 7.83 4.14 ;
      RECT 6.63 2.035 7.73 2.265 ;
      RECT 7.215 2.54 7.5 3.11 ;
      RECT 7.16 2.54 7.215 3 ;
      RECT 6.515 2.76 7.16 3 ;
      RECT 6.895 1.085 7.125 1.745 ;
      RECT 6.64 1.085 6.895 1.315 ;
      RECT 6.575 2.035 6.63 2.4 ;
      RECT 6.345 1.6 6.575 2.4 ;
      RECT 6.285 2.76 6.515 4.225 ;
      RECT 5.745 1.6 6.345 1.83 ;
      RECT 6.29 2.06 6.345 2.4 ;
      RECT 6.055 2.76 6.285 2.99 ;
      RECT 2.43 3.995 6.285 4.225 ;
      RECT 5.96 2.225 6.055 2.99 ;
      RECT 5.825 2.115 5.96 2.99 ;
      RECT 5.62 2.115 5.825 2.455 ;
      RECT 5.515 0.63 5.745 1.83 ;
      RECT 5.59 3.315 5.72 3.655 ;
      RECT 5.38 2.705 5.59 3.655 ;
      RECT 4.43 0.63 5.515 0.86 ;
      RECT 5.36 2.705 5.38 3.6 ;
      RECT 5.085 2.705 5.36 2.935 ;
      RECT 5.085 1.13 5.285 1.69 ;
      RECT 5.055 1.13 5.085 2.935 ;
      RECT 4.855 1.46 5.055 2.935 ;
      RECT 4.525 3.32 4.865 3.66 ;
      RECT 4.745 1.905 4.855 2.245 ;
      RECT 4.515 1.145 4.54 1.485 ;
      RECT 4.52 3.32 4.525 3.605 ;
      RECT 4.515 2.625 4.52 3.605 ;
      RECT 4.43 1.145 4.515 3.605 ;
      RECT 4.29 0.63 4.43 3.605 ;
      RECT 4.285 0.63 4.29 3.55 ;
      RECT 4.2 0.63 4.285 1.485 ;
      RECT 3.86 2.625 4.285 2.855 ;
      RECT 4 1.945 4.055 2.175 ;
      RECT 3.77 1.94 4 2.175 ;
      RECT 3.52 2.57 3.86 2.91 ;
      RECT 2.89 1.94 3.77 2.17 ;
      RECT 2.66 1.115 2.89 3.59 ;
      RECT 2.12 1.115 2.66 1.345 ;
      RECT 2.2 1.96 2.43 4.225 ;
      RECT 2.1 1.96 2.2 2.19 ;
      RECT 0.61 3.995 2.2 4.225 ;
      RECT 1.87 1.695 2.1 2.19 ;
      RECT 0.39 2.89 0.61 4.225 ;
      RECT 0.39 1.445 0.54 1.785 ;
      RECT 0.38 1.445 0.39 4.225 ;
      RECT 0.27 1.445 0.38 4.19 ;
      RECT 0.2 1.445 0.27 3.12 ;
      RECT 0.16 1.55 0.2 3.12 ;
  END
END DFFHQX4

MACRO DFFHQX2
  CLASS CORE ;
  FOREIGN DFFHQX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.2 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFHQXL ;

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8394 ;
  ANTENNAPARTIALMETALAREA 0.8163 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9008 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.9 0.7 12.24 1.04 ;
      RECT 11.525 0.81 11.9 1.04 ;
      RECT 11.525 2.94 11.74 3.22 ;
      RECT 11.295 0.81 11.525 3.22 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.144 ;
  ANTENNAPARTIALMETALAREA 0.335 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.325 1.405 1.825 2.075 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2628 ;
  ANTENNAPARTIALMETALAREA 0.2691 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1448 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.38 1.49 2.77 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13 -0.4 13.2 0.4 ;
      RECT 12.66 -0.4 13 0.95 ;
      RECT 11.44 -0.4 12.66 0.4 ;
      RECT 11.1 -0.4 11.44 0.575 ;
      RECT 9.425 -0.4 11.1 0.4 ;
      RECT 9.195 -0.4 9.425 1.075 ;
      RECT 6.32 -0.4 9.195 0.4 ;
      RECT 5.98 -0.4 6.32 1.44 ;
      RECT 4.02 -0.4 5.98 0.4 ;
      RECT 3.68 -0.4 4.02 1.27 ;
      RECT 1.08 -0.4 3.68 0.4 ;
      RECT 0.74 -0.4 1.08 0.575 ;
      RECT 0 -0.4 0.74 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.34 4.64 13.2 5.44 ;
      RECT 12 4.465 12.34 5.44 ;
      RECT 10.36 4.64 12 5.44 ;
      RECT 8.61 4.465 10.36 5.44 ;
      RECT 5.91 4.64 8.61 5.44 ;
      RECT 5.57 4.465 5.91 5.44 ;
      RECT 1.97 4.64 5.57 5.44 ;
      RECT 1.63 4.465 1.97 5.44 ;
      RECT 0 4.64 1.63 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.435 1.515 12.665 4.14 ;
      RECT 11.9 1.515 12.435 1.745 ;
      RECT 11.58 3.91 12.435 4.14 ;
      RECT 11.97 2.285 12.2 3.68 ;
      RECT 11.065 3.45 11.97 3.68 ;
      RECT 11.235 3.91 11.58 4.37 ;
      RECT 10.605 3.91 11.235 4.14 ;
      RECT 10.835 1.5 11.065 3.68 ;
      RECT 10.28 1.5 10.835 1.73 ;
      RECT 9.45 3.36 10.835 3.59 ;
      RECT 10.375 1.96 10.605 3.13 ;
      RECT 10.375 3.905 10.605 4.14 ;
      RECT 8.465 1.96 10.375 2.19 ;
      RECT 8.195 2.9 10.375 3.13 ;
      RECT 10.06 3.905 10.375 4.135 ;
      RECT 9.94 1.165 10.28 1.73 ;
      RECT 7.47 2.42 10.07 2.65 ;
      RECT 8.925 1.5 9.94 1.73 ;
      RECT 9.34 3.36 9.45 3.7 ;
      RECT 9.11 3.36 9.34 4.135 ;
      RECT 7.13 3.905 9.11 4.135 ;
      RECT 8.695 0.64 8.925 1.73 ;
      RECT 7.95 0.64 8.695 0.87 ;
      RECT 8.235 1.1 8.465 2.19 ;
      RECT 7.025 1.445 8.235 1.675 ;
      RECT 7.965 2.9 8.195 3.675 ;
      RECT 7.85 3.39 7.965 3.675 ;
      RECT 7.72 0.64 7.95 1.215 ;
      RECT 6.695 3.39 7.85 3.62 ;
      RECT 7.46 0.985 7.72 1.215 ;
      RECT 7.36 2.42 7.47 3.16 ;
      RECT 7.13 1.905 7.36 3.16 ;
      RECT 5.51 1.905 7.13 2.135 ;
      RECT 6.235 2.93 7.13 3.16 ;
      RECT 6.795 1.1 7.025 1.675 ;
      RECT 6.465 3.39 6.695 3.73 ;
      RECT 5.775 2.365 6.61 2.595 ;
      RECT 6.005 2.93 6.235 4.235 ;
      RECT 2.375 4.005 6.005 4.235 ;
      RECT 5.545 2.365 5.775 3.775 ;
      RECT 4.765 3.545 5.545 3.775 ;
      RECT 5.375 1.105 5.52 1.445 ;
      RECT 5.28 0.63 5.375 1.445 ;
      RECT 5.28 2.365 5.315 2.965 ;
      RECT 5.085 0.63 5.28 2.965 ;
      RECT 5.05 0.63 5.085 2.595 ;
      RECT 5.015 0.63 5.05 0.86 ;
      RECT 4.535 0.95 4.765 3.775 ;
      RECT 3.625 2.16 4.535 2.5 ;
      RECT 3.395 1.545 4.18 1.775 ;
      RECT 3.165 1.545 3.395 3.6 ;
      RECT 2.97 1.545 3.165 1.775 ;
      RECT 2.74 0.92 2.97 1.775 ;
      RECT 2.66 0.92 2.74 1.15 ;
      RECT 2.32 0.81 2.66 1.15 ;
      RECT 2.375 1.38 2.43 1.72 ;
      RECT 2.145 1.38 2.375 4.235 ;
      RECT 2.09 1.38 2.145 1.72 ;
      RECT 1.21 3.135 2.145 3.365 ;
      RECT 0.87 3.025 1.21 3.365 ;
      RECT 0.57 3.025 0.87 3.255 ;
      RECT 0.34 1.34 0.57 3.255 ;
      RECT 0.18 1.34 0.34 1.68 ;
  END
END DFFHQX2

MACRO DFFHQX1
  CLASS CORE ;
  FOREIGN DFFHQX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFHQXL ;

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5176 ;
  ANTENNAPARTIALMETALAREA 1.2379 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.3636 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.345 0.695 10.435 3.53 ;
      RECT 10.205 0.695 10.345 3.755 ;
      RECT 9.59 0.695 10.205 0.925 ;
      RECT 10.115 3.19 10.205 3.755 ;
      RECT 9.05 3.19 10.115 3.53 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3483 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3144 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.41 1.82 1.84 2.63 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2016 ;
  ANTENNAPARTIALMETALAREA 0.256 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.205 1.18 2.66 ;
      RECT 0.645 2.15 0.875 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.17 -0.4 10.56 0.4 ;
      RECT 8.83 -0.4 9.17 0.575 ;
      RECT 6.315 -0.4 8.83 0.4 ;
      RECT 6.085 -0.4 6.315 1.46 ;
      RECT 4.015 -0.4 6.085 0.4 ;
      RECT 3.785 -0.4 4.015 1.15 ;
      RECT 1.35 -0.4 3.785 0.4 ;
      RECT 1.01 -0.4 1.35 0.575 ;
      RECT 0 -0.4 1.01 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.12 4.64 10.56 5.44 ;
      RECT 9.78 4.41 10.12 5.44 ;
      RECT 8.63 4.64 9.78 5.44 ;
      RECT 8.29 4.465 8.63 5.44 ;
      RECT 5.795 4.64 8.29 5.44 ;
      RECT 5.455 4.465 5.795 5.44 ;
      RECT 1.815 4.64 5.455 5.44 ;
      RECT 1.475 4.465 1.815 5.44 ;
      RECT 0 4.64 1.475 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.925 1.46 9.97 1.8 ;
      RECT 9.695 1.46 9.925 2.96 ;
      RECT 9.63 1.46 9.695 1.8 ;
      RECT 8.64 2.73 9.695 2.96 ;
      RECT 9.235 2.04 9.465 2.38 ;
      RECT 9.09 4.115 9.39 4.345 ;
      RECT 9.17 2.04 9.235 2.27 ;
      RECT 8.94 1.605 9.17 2.27 ;
      RECT 8.86 4.005 9.09 4.345 ;
      RECT 7.955 1.605 8.94 1.835 ;
      RECT 8.64 4.005 8.86 4.235 ;
      RECT 8.41 2.18 8.64 4.235 ;
      RECT 8.3 2.18 8.41 2.52 ;
      RECT 6.775 0.875 8.39 1.105 ;
      RECT 7.725 1.44 7.955 4.375 ;
      RECT 7.03 4.145 7.725 4.375 ;
      RECT 7.265 1.445 7.495 3.915 ;
      RECT 7.235 1.445 7.265 1.675 ;
      RECT 6.595 3.685 7.265 3.915 ;
      RECT 7.005 1.335 7.235 1.675 ;
      RECT 6.865 2.82 7.035 3.165 ;
      RECT 6.775 1.905 6.865 3.455 ;
      RECT 6.635 0.875 6.775 3.455 ;
      RECT 6.545 0.875 6.635 2.135 ;
      RECT 6.135 3.225 6.635 3.455 ;
      RECT 6.365 3.685 6.595 4.185 ;
      RECT 5.905 1.905 6.545 2.135 ;
      RECT 6.135 2.38 6.365 2.995 ;
      RECT 5.675 2.765 6.135 2.995 ;
      RECT 5.905 3.225 6.135 4.235 ;
      RECT 5.675 1.765 5.905 2.135 ;
      RECT 2.375 4.005 5.905 4.235 ;
      RECT 5.56 1.765 5.675 1.995 ;
      RECT 5.445 2.765 5.675 3.775 ;
      RECT 5.365 1.17 5.57 1.51 ;
      RECT 4.625 3.545 5.445 3.775 ;
      RECT 5.275 0.63 5.365 1.51 ;
      RECT 5.215 0.63 5.275 1.615 ;
      RECT 5.135 0.63 5.215 3.13 ;
      RECT 5.045 1.225 5.135 3.13 ;
      RECT 4.985 1.385 5.045 3.13 ;
      RECT 4.625 0.81 4.815 1.155 ;
      RECT 4.585 0.81 4.625 3.775 ;
      RECT 4.395 0.925 4.585 3.775 ;
      RECT 3.92 2.185 4.395 2.415 ;
      RECT 3.935 1.455 4.165 1.8 ;
      RECT 3.295 1.455 3.935 1.685 ;
      RECT 3.58 2.13 3.92 2.47 ;
      RECT 3.065 0.805 3.295 3.68 ;
      RECT 2.37 0.805 3.065 1.035 ;
      RECT 2.145 1.39 2.375 4.235 ;
      RECT 1.055 3.135 2.145 3.365 ;
      RECT 0.715 3.025 1.055 3.365 ;
      RECT 0.415 1.43 0.75 1.77 ;
      RECT 0.415 3.025 0.715 3.255 ;
      RECT 0.41 1.43 0.415 3.255 ;
      RECT 0.185 1.54 0.41 3.255 ;
  END
END DFFHQX1

MACRO DFFXL
  CLASS CORE ;
  FOREIGN DFFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.22 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6466 ;
  ANTENNAPARTIALMETALAREA 0.8479 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.0227 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.345 3.515 10.435 3.855 ;
      RECT 10.28 0.81 10.345 3.855 ;
      RECT 10.115 0.705 10.28 3.855 ;
      RECT 10.05 0.705 10.115 1.285 ;
      RECT 10.095 3.515 10.115 3.855 ;
      RECT 9.81 0.705 10.05 0.935 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.442 ;
  ANTENNAPARTIALMETALAREA 1.085 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.1887 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.18 0.685 9.45 0.915 ;
      RECT 9.115 1.875 9.345 3.44 ;
      RECT 9.01 0.685 9.18 1.165 ;
      RECT 9.01 1.875 9.115 2.105 ;
      RECT 9.075 3.21 9.115 3.44 ;
      RECT 8.735 3.21 9.075 3.55 ;
      RECT 8.95 0.685 9.01 2.105 ;
      RECT 8.78 0.935 8.95 2.105 ;
      RECT 8.135 1.285 8.78 1.515 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.635 1.845 1.765 2.075 ;
      RECT 1.35 1.475 1.635 2.075 ;
      RECT 1.295 1.475 1.35 1.815 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2133 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.305 1.18 2.66 ;
      RECT 0.8 2.2 0.875 2.66 ;
      RECT 0.645 2.2 0.8 2.655 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.85 -0.4 11.22 0.4 ;
      RECT 10.51 -0.4 10.85 0.575 ;
      RECT 8.69 -0.4 10.51 0.4 ;
      RECT 8.35 -0.4 8.69 0.575 ;
      RECT 6.25 -0.4 8.35 0.4 ;
      RECT 5.91 -0.4 6.25 1.51 ;
      RECT 3.895 -0.4 5.91 0.4 ;
      RECT 3.665 -0.4 3.895 1.15 ;
      RECT 1.175 -0.4 3.665 0.4 ;
      RECT 0.835 -0.4 1.175 0.575 ;
      RECT 0 -0.4 0.835 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.735 4.64 11.22 5.44 ;
      RECT 9.395 4.41 9.735 5.44 ;
      RECT 8.275 4.64 9.395 5.44 ;
      RECT 7.935 4.465 8.275 5.44 ;
      RECT 5.795 4.64 7.935 5.44 ;
      RECT 5.455 4.465 5.795 5.44 ;
      RECT 1.38 4.64 5.455 5.44 ;
      RECT 1.04 4.41 1.38 5.44 ;
      RECT 0 4.64 1.04 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.58 1.415 9.81 4.18 ;
      RECT 9.24 1.415 9.58 1.645 ;
      RECT 9.095 3.95 9.58 4.18 ;
      RECT 8.865 3.95 9.095 4.35 ;
      RECT 8.645 4.005 8.865 4.35 ;
      RECT 8.31 2.67 8.795 2.9 ;
      RECT 7.85 4.005 8.645 4.235 ;
      RECT 8.08 2.26 8.31 2.9 ;
      RECT 7.53 2.26 8.08 2.49 ;
      RECT 6.775 0.67 7.93 0.9 ;
      RECT 7.62 2.745 7.85 4.235 ;
      RECT 7.24 1.27 7.53 2.49 ;
      RECT 7.19 1.27 7.24 4.15 ;
      RECT 7.115 2.26 7.19 4.15 ;
      RECT 7.01 2.26 7.115 4.26 ;
      RECT 6.775 3.92 7.01 4.26 ;
      RECT 6.665 0.67 6.775 3.26 ;
      RECT 6.545 0.67 6.665 3.615 ;
      RECT 5.665 1.74 6.545 1.97 ;
      RECT 6.435 2.92 6.545 3.615 ;
      RECT 6.27 3.385 6.435 3.615 ;
      RECT 6.205 2.2 6.31 2.69 ;
      RECT 6.04 3.385 6.27 4.235 ;
      RECT 6.08 2.2 6.205 3.135 ;
      RECT 5.975 2.46 6.08 3.135 ;
      RECT 2.79 4.005 6.04 4.235 ;
      RECT 5.8 2.905 5.975 3.135 ;
      RECT 5.57 2.905 5.8 3.775 ;
      RECT 5.59 1.74 5.665 2.325 ;
      RECT 5.435 1.74 5.59 2.51 ;
      RECT 4.66 3.545 5.57 3.775 ;
      RECT 5.245 1.17 5.45 1.51 ;
      RECT 5.36 2.095 5.435 2.51 ;
      RECT 5.175 0.63 5.245 1.51 ;
      RECT 5.13 2.78 5.235 3.12 ;
      RECT 5.13 0.63 5.175 1.61 ;
      RECT 5.015 0.63 5.13 3.12 ;
      RECT 4.945 1.225 5.015 3.12 ;
      RECT 4.9 1.38 4.945 3.12 ;
      RECT 4.895 2.78 4.9 3.12 ;
      RECT 4.66 0.81 4.695 1.15 ;
      RECT 4.465 0.81 4.66 3.775 ;
      RECT 4.43 0.92 4.465 3.775 ;
      RECT 3.865 2.455 4.43 2.685 ;
      RECT 3.375 1.785 4.2 2.015 ;
      RECT 3.525 2.4 3.865 2.74 ;
      RECT 3.25 0.795 3.375 2.015 ;
      RECT 3.02 0.795 3.25 3.68 ;
      RECT 2.25 0.795 3.02 1.025 ;
      RECT 2.56 3.25 2.79 4.235 ;
      RECT 2.315 3.25 2.56 3.48 ;
      RECT 2.085 1.39 2.315 3.48 ;
      RECT 0.54 3.25 2.085 3.48 ;
      RECT 0.38 3.14 0.54 3.48 ;
      RECT 0.38 1.065 0.52 1.405 ;
      RECT 0.2 1.065 0.38 3.48 ;
      RECT 0.18 1.065 0.2 3.37 ;
      RECT 0.15 1.12 0.18 3.37 ;
  END
END DFFXL

MACRO DFFX4
  CLASS CORE ;
  FOREIGN DFFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 16.5 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5876 ;
  ANTENNAPARTIALMETALAREA 1.2674 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.3725 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.19 0.77 15.53 1.58 ;
      RECT 15.05 2.865 15.39 3.675 ;
      RECT 15.045 1.2 15.19 1.58 ;
      RECT 15.04 2.865 15.05 3.095 ;
      RECT 15.04 1.2 15.045 2.075 ;
      RECT 14.81 1.2 15.04 3.095 ;
      RECT 14.66 1.2 14.81 2.66 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5876 ;
  ANTENNAPARTIALMETALAREA 1.2488 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7206 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.89 0.835 14.01 1.645 ;
      RECT 13.87 0.835 13.89 3.385 ;
      RECT 13.67 0.835 13.87 3.675 ;
      RECT 13.66 1.125 13.67 3.675 ;
      RECT 13.53 1.82 13.66 3.675 ;
      RECT 13.34 1.82 13.53 3.22 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2988 ;
  ANTENNAPARTIALMETALAREA 0.3096 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5953 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.745 2.405 1.765 2.635 ;
      RECT 1.74 1.55 1.745 2.635 ;
      RECT 1.51 1.495 1.74 2.635 ;
      RECT 1.4 1.495 1.51 1.835 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.4788 ;
  ANTENNAPARTIALMETALAREA 0.2283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.58 2.2 1.105 2.635 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.31 -0.4 16.5 0.4 ;
      RECT 15.97 -0.4 16.31 0.575 ;
      RECT 14.77 -0.4 15.97 0.4 ;
      RECT 14.43 -0.4 14.77 0.575 ;
      RECT 13.235 -0.4 14.43 0.4 ;
      RECT 13.005 -0.4 13.235 1.35 ;
      RECT 11.795 -0.4 13.005 0.4 ;
      RECT 11.565 -0.4 11.795 1.31 ;
      RECT 9.155 -0.4 11.565 0.4 ;
      RECT 8.925 -0.4 9.155 1.335 ;
      RECT 6.595 -0.4 8.925 0.4 ;
      RECT 6.365 -0.4 6.595 1.37 ;
      RECT 4.1 -0.4 6.365 0.4 ;
      RECT 3.76 -0.4 4.1 1.27 ;
      RECT 1.365 -0.4 3.76 0.4 ;
      RECT 1.025 -0.4 1.365 0.575 ;
      RECT 0 -0.4 1.025 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.15 4.64 16.5 5.44 ;
      RECT 15.81 4.465 16.15 5.44 ;
      RECT 14.63 4.64 15.81 5.44 ;
      RECT 14.29 4.465 14.63 5.44 ;
      RECT 13.11 4.64 14.29 5.44 ;
      RECT 12.77 4.465 13.11 5.44 ;
      RECT 11.79 4.64 12.77 5.44 ;
      RECT 11.45 4.465 11.79 5.44 ;
      RECT 9.345 4.64 11.45 5.44 ;
      RECT 9.005 4.005 9.345 5.44 ;
      RECT 6.52 4.64 9.005 5.44 ;
      RECT 6.18 4.465 6.52 5.44 ;
      RECT 3.03 4.64 6.18 5.44 ;
      RECT 2.575 4.465 3.03 5.44 ;
      RECT 1.38 4.64 2.575 5.44 ;
      RECT 1.04 4.465 1.38 5.44 ;
      RECT 0 4.64 1.04 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.715 2.33 15.945 4.16 ;
      RECT 15.62 2.33 15.715 2.56 ;
      RECT 13.095 3.93 15.715 4.16 ;
      RECT 15.39 2.055 15.62 2.56 ;
      RECT 12.865 2.115 13.095 4.16 ;
      RECT 12.515 2.115 12.865 2.345 ;
      RECT 12.21 3.47 12.865 3.81 ;
      RECT 12.285 1.04 12.515 2.345 ;
      RECT 11.325 2.785 12.49 3.015 ;
      RECT 11.6 2.115 12.285 2.345 ;
      RECT 11.095 0.97 11.325 3.49 ;
      RECT 10.49 0.97 11.095 1.25 ;
      RECT 10.63 3.26 11.095 3.49 ;
      RECT 10.26 1.55 10.86 1.78 ;
      RECT 10.29 3.26 10.63 4.07 ;
      RECT 10.15 0.965 10.49 1.305 ;
      RECT 8.06 3.45 10.29 3.68 ;
      RECT 10.205 1.55 10.26 2.935 ;
      RECT 10.03 1.55 10.205 2.97 ;
      RECT 9.8 1.075 10.15 1.305 ;
      RECT 9.92 2.595 10.03 2.97 ;
      RECT 9.755 2.74 9.92 2.97 ;
      RECT 9.57 1.075 9.8 1.805 ;
      RECT 9.525 2.74 9.755 3.04 ;
      RECT 8.53 1.575 9.57 1.805 ;
      RECT 8.3 2.81 9.525 3.04 ;
      RECT 9.23 2.235 9.285 2.575 ;
      RECT 8.945 2.035 9.23 2.575 ;
      RECT 7.02 2.035 8.945 2.265 ;
      RECT 8.3 1.25 8.53 1.805 ;
      RECT 7.93 1.25 8.3 1.48 ;
      RECT 8.015 2.595 8.3 3.04 ;
      RECT 7.72 3.45 8.06 4.26 ;
      RECT 7.96 2.595 8.015 3 ;
      RECT 6.795 2.76 7.96 3 ;
      RECT 7.59 1.14 7.93 1.48 ;
      RECT 6.965 2.035 7.02 2.4 ;
      RECT 6.735 1.6 6.965 2.4 ;
      RECT 6.565 2.76 6.795 4.225 ;
      RECT 6.135 1.6 6.735 1.83 ;
      RECT 6.68 2.06 6.735 2.4 ;
      RECT 6.445 2.76 6.565 2.99 ;
      RECT 3.535 3.995 6.565 4.225 ;
      RECT 6.35 2.225 6.445 2.99 ;
      RECT 6.215 2.115 6.35 2.99 ;
      RECT 6.01 2.115 6.215 2.455 ;
      RECT 5.905 0.63 6.135 1.83 ;
      RECT 5.98 3.315 6.11 3.655 ;
      RECT 5.77 2.705 5.98 3.655 ;
      RECT 4.82 0.63 5.905 0.86 ;
      RECT 5.75 2.705 5.77 3.6 ;
      RECT 5.31 2.705 5.75 2.935 ;
      RECT 5.445 1.175 5.675 1.69 ;
      RECT 5.37 1.46 5.445 1.69 ;
      RECT 5.365 1.46 5.37 2.19 ;
      RECT 5.31 1.46 5.365 2.245 ;
      RECT 5.14 1.46 5.31 2.935 ;
      RECT 4.805 3.32 5.145 3.66 ;
      RECT 5.08 1.905 5.14 2.935 ;
      RECT 5.025 1.905 5.08 2.245 ;
      RECT 4.795 0.63 4.82 1.485 ;
      RECT 4.8 3.32 4.805 3.605 ;
      RECT 4.795 2.625 4.8 3.605 ;
      RECT 4.59 0.63 4.795 3.605 ;
      RECT 4.57 1.145 4.59 3.605 ;
      RECT 4.565 1.145 4.57 3.55 ;
      RECT 4.48 1.145 4.565 1.485 ;
      RECT 4.14 2.625 4.565 2.855 ;
      RECT 4.28 1.945 4.335 2.175 ;
      RECT 4.05 1.94 4.28 2.175 ;
      RECT 3.8 2.57 4.14 2.91 ;
      RECT 3.17 1.94 4.05 2.17 ;
      RECT 3.25 3.89 3.535 4.225 ;
      RECT 2.71 3.89 3.25 4.15 ;
      RECT 2.94 0.685 3.17 3.59 ;
      RECT 2.4 0.685 2.94 0.915 ;
      RECT 2.48 2.82 2.71 4.15 ;
      RECT 2.36 2.82 2.48 3.05 ;
      RECT 1.84 3.92 2.48 4.15 ;
      RECT 2.13 1.39 2.36 3.05 ;
      RECT 1.61 3.92 1.84 4.235 ;
      RECT 0.62 4.005 1.61 4.235 ;
      RECT 0.35 2.87 0.62 4.235 ;
      RECT 0.35 0.845 0.52 1.655 ;
      RECT 0.28 0.845 0.35 4.235 ;
      RECT 0.18 0.845 0.28 3.255 ;
      RECT 0.12 1.135 0.18 3.255 ;
  END
END DFFX4

MACRO DFFX2
  CLASS CORE ;
  FOREIGN DFFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.81 ;
  ANTENNAPARTIALMETALAREA 0.6532 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0581 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.755 1.355 12.985 3.33 ;
      RECT 12.68 1.355 12.755 1.845 ;
      RECT 12.7 3.1 12.755 3.33 ;
      RECT 12.36 3.1 12.7 3.44 ;
      RECT 12.58 1.355 12.68 1.695 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.858 ;
  ANTENNAPARTIALMETALAREA 0.852 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9538 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.505 0.7 11.56 1.04 ;
      RECT 11.22 0.7 11.505 1.08 ;
      RECT 10.865 0.85 11.22 1.08 ;
      RECT 11.08 2.87 11.16 3.21 ;
      RECT 10.865 2.38 11.08 3.21 ;
      RECT 10.82 0.85 10.865 3.21 ;
      RECT 10.7 0.85 10.82 2.66 ;
      RECT 10.635 0.85 10.7 2.61 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.162 ;
  ANTENNAPARTIALMETALAREA 0.2904 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.405 1.825 2.075 ;
      RECT 1.325 1.405 1.46 1.745 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2052 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9752 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.12 1.18 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.48 -0.4 13.86 0.4 ;
      RECT 13.14 -0.4 13.48 0.575 ;
      RECT 12.36 -0.4 13.14 0.4 ;
      RECT 12.02 -0.4 12.36 0.575 ;
      RECT 10.76 -0.4 12.02 0.4 ;
      RECT 10.42 -0.4 10.76 0.575 ;
      RECT 8.8 -0.4 10.42 0.4 ;
      RECT 8.46 -0.4 8.8 1.27 ;
      RECT 6.185 -0.4 8.46 0.4 ;
      RECT 5.845 -0.4 6.185 1.445 ;
      RECT 4.02 -0.4 5.845 0.4 ;
      RECT 3.68 -0.4 4.02 1.27 ;
      RECT 1.1 -0.4 3.68 0.4 ;
      RECT 0.76 -0.4 1.1 0.575 ;
      RECT 0 -0.4 0.76 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.26 4.64 13.86 5.44 ;
      RECT 12.92 4.465 13.26 5.44 ;
      RECT 11.92 4.64 12.92 5.44 ;
      RECT 11.58 4.465 11.92 5.44 ;
      RECT 9.94 4.64 11.58 5.44 ;
      RECT 8.19 4.465 9.94 5.44 ;
      RECT 5.89 4.64 8.19 5.44 ;
      RECT 5.55 4.465 5.89 5.44 ;
      RECT 4.53 4.64 5.55 5.44 ;
      RECT 4.19 4.465 4.53 5.44 ;
      RECT 1.45 4.64 4.19 5.44 ;
      RECT 1.11 4.41 1.45 5.44 ;
      RECT 0 4.64 1.11 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.435 4.02 12.49 4.36 ;
      RECT 12.15 3.995 12.435 4.36 ;
      RECT 12.125 3.995 12.15 4.225 ;
      RECT 11.895 1.545 12.125 4.225 ;
      RECT 11.22 1.545 11.895 1.775 ;
      RECT 11.16 3.995 11.895 4.225 ;
      RECT 11.435 2.285 11.665 3.67 ;
      RECT 9.975 3.44 11.435 3.67 ;
      RECT 11.05 3.995 11.16 4.37 ;
      RECT 10.82 3.9 11.05 4.37 ;
      RECT 9.64 3.9 10.82 4.13 ;
      RECT 9.745 1.775 9.975 3.67 ;
      RECT 9.6 1.775 9.745 2.005 ;
      RECT 9.03 3.36 9.745 3.67 ;
      RECT 9.37 1.155 9.6 2.005 ;
      RECT 9.11 2.35 9.45 2.69 ;
      RECT 9.26 1.155 9.37 1.795 ;
      RECT 8.13 1.565 9.26 1.795 ;
      RECT 8.195 2.405 9.11 2.635 ;
      RECT 8.92 3.36 9.03 3.7 ;
      RECT 8.69 3.36 8.92 3.96 ;
      RECT 7.155 3.73 8.69 3.96 ;
      RECT 7.965 2.405 8.195 3.16 ;
      RECT 7.9 1.16 8.13 1.795 ;
      RECT 7.3 2.93 7.965 3.16 ;
      RECT 7.52 1.16 7.9 1.39 ;
      RECT 7.18 1.05 7.52 1.39 ;
      RECT 7.21 2.82 7.3 3.16 ;
      RECT 6.98 1.785 7.21 3.16 ;
      RECT 6.925 3.44 7.155 4.275 ;
      RECT 5.53 1.785 6.98 2.015 ;
      RECT 6.96 2.82 6.98 3.16 ;
      RECT 6.33 2.93 6.96 3.16 ;
      RECT 5.86 2.245 6.61 2.475 ;
      RECT 6.1 2.93 6.33 4.235 ;
      RECT 3.595 4.005 6.1 4.235 ;
      RECT 5.63 2.245 5.86 3.775 ;
      RECT 4.695 3.545 5.63 3.775 ;
      RECT 5.295 1.105 5.445 1.445 ;
      RECT 5.295 2.625 5.33 2.965 ;
      RECT 5.065 0.63 5.295 2.965 ;
      RECT 4.935 0.63 5.065 0.86 ;
      RECT 4.99 2.625 5.065 2.965 ;
      RECT 4.685 2.27 4.695 3.775 ;
      RECT 4.465 0.95 4.685 3.775 ;
      RECT 4.455 0.95 4.465 2.51 ;
      RECT 3.585 2.17 4.455 2.51 ;
      RECT 3.355 1.555 4.18 1.785 ;
      RECT 3.365 3.89 3.595 4.235 ;
      RECT 3.31 3.89 3.365 4.225 ;
      RECT 3.125 1.545 3.355 3.6 ;
      RECT 3.3 3.89 3.31 4.15 ;
      RECT 2.895 3.89 3.3 4.12 ;
      RECT 2.97 1.545 3.125 1.785 ;
      RECT 2.74 0.92 2.97 1.785 ;
      RECT 2.665 2.82 2.895 4.12 ;
      RECT 2.66 0.92 2.74 1.15 ;
      RECT 2.375 2.82 2.665 3.05 ;
      RECT 1.98 3.89 2.665 4.12 ;
      RECT 2.32 0.81 2.66 1.15 ;
      RECT 2.375 1.38 2.43 1.72 ;
      RECT 2.145 1.38 2.375 3.05 ;
      RECT 2.09 1.38 2.145 1.72 ;
      RECT 1.75 3.605 1.98 4.12 ;
      RECT 1.31 3.605 1.75 3.835 ;
      RECT 0.91 3.02 1.31 3.835 ;
      RECT 0.57 3.08 0.91 3.31 ;
      RECT 0.34 1.34 0.57 3.31 ;
      RECT 0.18 1.34 0.34 1.68 ;
  END
END DFFX2

MACRO DFFX1
  CLASS CORE ;
  FOREIGN DFFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.22 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ DFFXL ;

  PIN QN
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.936 ;
  ANTENNAPARTIALMETALAREA 0.9486 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3178 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.7 1.19 11.04 3.88 ;
      RECT 10.6 3.54 10.7 3.88 ;
     END
  END QN

  PIN Q
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.532 ;
  ANTENNAPARTIALMETALAREA 1.1843 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.115 0.865 10.345 3.42 ;
      RECT 9.83 0.865 10.115 1.095 ;
      RECT 9.23 3.19 10.115 3.42 ;
      RECT 9.3 0.695 9.83 1.095 ;
      RECT 8.89 3.19 9.23 3.53 ;
     END
  END Q

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2456 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2137 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.69 1.845 1.765 2.075 ;
      RECT 1.41 1.405 1.69 2.075 ;
      RECT 1.29 1.405 1.41 1.745 ;
     END
  END D

  PIN CK
  DIRECTION INPUT ;
  USE CLOCK ;
  ANTENNAGATEAREA 0.1908 ;
  ANTENNAPARTIALMETALAREA 0.2265 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.94 2.205 1.18 2.66 ;
      RECT 0.71 2.15 0.94 2.66 ;
     END
  END CK

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.46 -0.4 11.22 0.4 ;
      RECT 10.12 -0.4 10.46 0.575 ;
      RECT 8.88 -0.4 10.12 0.4 ;
      RECT 8.54 -0.4 8.88 0.575 ;
      RECT 6.44 -0.4 8.54 0.4 ;
      RECT 6.1 -0.4 6.44 1.46 ;
      RECT 4.015 -0.4 6.1 0.4 ;
      RECT 3.785 -0.4 4.015 1.15 ;
      RECT 1.225 -0.4 3.785 0.4 ;
      RECT 0.885 -0.4 1.225 0.575 ;
      RECT 0 -0.4 0.885 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.18 4.64 11.22 5.44 ;
      RECT 9.84 4.41 10.18 5.44 ;
      RECT 8.47 4.64 9.84 5.44 ;
      RECT 8.13 4.465 8.47 5.44 ;
      RECT 5.795 4.64 8.13 5.44 ;
      RECT 5.455 4.465 5.795 5.44 ;
      RECT 1.55 4.64 5.455 5.44 ;
      RECT 1.21 4.465 1.55 5.44 ;
      RECT 0 4.64 1.21 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 9.68 1.6 9.87 2.765 ;
      RECT 9.64 1.49 9.68 2.765 ;
      RECT 9.34 1.49 9.64 1.83 ;
      RECT 8.4 2.535 9.64 2.765 ;
      RECT 8.88 2.075 9.255 2.305 ;
      RECT 9.11 4.14 9.23 4.37 ;
      RECT 8.88 3.97 9.11 4.37 ;
      RECT 8.65 1.44 8.88 2.305 ;
      RECT 8.4 3.97 8.88 4.2 ;
      RECT 7.55 1.44 8.65 1.835 ;
      RECT 8.35 2.535 8.4 4.2 ;
      RECT 8.17 2.18 8.35 4.2 ;
      RECT 8.12 2.18 8.17 2.765 ;
      RECT 8.01 2.18 8.12 2.52 ;
      RECT 6.94 0.875 8.1 1.105 ;
      RECT 7.32 1.44 7.55 4.285 ;
      RECT 6.87 4.055 7.32 4.285 ;
      RECT 6.94 2.82 7.09 3.16 ;
      RECT 6.865 0.875 6.94 3.16 ;
      RECT 6.71 0.875 6.865 3.615 ;
      RECT 6.635 1.765 6.71 3.615 ;
      RECT 5.56 1.765 6.635 1.995 ;
      RECT 6.27 3.385 6.635 3.615 ;
      RECT 6.135 2.38 6.365 3.135 ;
      RECT 6.04 3.385 6.27 4.235 ;
      RECT 5.8 2.905 6.135 3.135 ;
      RECT 3.535 4.005 6.04 4.235 ;
      RECT 5.57 2.905 5.8 3.775 ;
      RECT 5.405 1.17 5.61 1.51 ;
      RECT 4.76 3.545 5.57 3.775 ;
      RECT 5.315 0.63 5.405 1.51 ;
      RECT 5.315 2.79 5.33 3.13 ;
      RECT 5.085 0.63 5.315 3.13 ;
      RECT 4.99 2.79 5.085 3.13 ;
      RECT 4.76 0.81 4.815 2.47 ;
      RECT 4.585 0.81 4.76 3.775 ;
      RECT 4.49 2.13 4.585 3.775 ;
      RECT 3.58 2.13 4.49 2.47 ;
      RECT 3.375 1.515 4.355 1.745 ;
      RECT 2.835 3.995 3.535 4.235 ;
      RECT 3.295 0.805 3.375 1.745 ;
      RECT 3.065 0.805 3.295 3.68 ;
      RECT 2.37 0.805 3.065 1.035 ;
      RECT 2.605 2.82 2.835 4.235 ;
      RECT 2.375 2.82 2.605 3.05 ;
      RECT 0.785 3.605 2.605 3.835 ;
      RECT 2.145 1.39 2.375 3.05 ;
      RECT 0.445 3.02 0.785 3.835 ;
      RECT 0.445 1.43 0.52 1.77 ;
      RECT 0.365 1.43 0.445 3.835 ;
      RECT 0.215 1.43 0.365 3.31 ;
      RECT 0.18 1.43 0.215 1.77 ;
  END
END DFFX1

MACRO CLKINVXL
  CLASS CORE ;
  FOREIGN CLKINVXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.98 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8008 ;
  ANTENNAPARTIALMETALAREA 1.1335 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4397 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.485 1.82 1.83 3.22 ;
      RECT 1.255 1.35 1.485 3.885 ;
      RECT 1.12 1.35 1.255 1.85 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1764 ;
  ANTENNAPARTIALMETALAREA 0.316 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.19 2.38 0.925 2.81 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 -0.4 1.98 0.4 ;
      RECT 0.98 -0.4 1.32 0.575 ;
      RECT 0 -0.4 0.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.89 4.64 1.98 5.44 ;
      RECT 0.525 4.395 0.89 5.44 ;
      RECT 0 4.64 0.525 5.44 ;
     END
  END VDD
END CLKINVXL

MACRO CLKINVX8
  CLASS CORE ;
  FOREIGN CLKINVX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.8133 ;
  ANTENNAPARTIALMETALAREA 4.122 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.8529 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.16 1.82 3.745 3.22 ;
      RECT 3.085 1.51 3.16 3.22 ;
      RECT 2.88 1.51 3.085 3.275 ;
      RECT 2.195 1.235 2.88 3.41 ;
      RECT 2.12 1.235 2.195 1.82 ;
      RECT 0.78 2.93 2.195 3.41 ;
      RECT 0.87 1.235 2.12 1.715 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.857 ;
  ANTENNAPARTIALMETALAREA 0.5012 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5158 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.54 2.045 1.355 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.005 -0.4 3.96 0.4 ;
      RECT 1.665 -0.4 2.005 0.98 ;
      RECT 0.56 -0.4 1.665 0.4 ;
      RECT 0.22 -0.4 0.56 0.575 ;
      RECT 0 -0.4 0.22 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.32 4.64 3.96 5.44 ;
      RECT 2.98 3.79 3.32 5.44 ;
      RECT 1.915 4.64 2.98 5.44 ;
      RECT 1.575 3.79 1.915 5.44 ;
      RECT 0.52 4.64 1.575 5.44 ;
      RECT 0.18 3.79 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
END CLKINVX8

MACRO CLKINVX4
  CLASS CORE ;
  FOREIGN CLKINVX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.323 ;
  ANTENNAPARTIALMETALAREA 1.5285 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.2771 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.29 1.84 3.78 ;
      RECT 1.08 1.29 1.46 1.67 ;
      RECT 1.44 2.965 1.46 3.78 ;
      RECT 1.1 2.965 1.44 4.205 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.882 ;
  ANTENNAPARTIALMETALAREA 0.5184 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.537 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.02 0.95 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.44 -0.4 2.64 0.4 ;
      RECT 2.1 -0.4 2.44 0.575 ;
      RECT 0.68 -0.4 2.1 0.4 ;
      RECT 0.34 -0.4 0.68 0.575 ;
      RECT 0 -0.4 0.34 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.2 4.64 2.64 5.44 ;
      RECT 1.86 4.465 2.2 5.44 ;
      RECT 0.68 4.64 1.86 5.44 ;
      RECT 0.34 4.465 0.68 5.44 ;
      RECT 0 4.64 0.34 5.44 ;
     END
  END VDD
END CLKINVX4

MACRO CLKINVX3
  CLASS CORE ;
  FOREIGN CLKINVX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.98 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.0164 ;
  ANTENNAPARTIALMETALAREA 0.7862 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9574 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.025 2.63 1.18 3.78 ;
      RECT 0.795 1.435 1.025 3.78 ;
      RECT 0.735 2.635 0.795 3.78 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6696 ;
  ANTENNAPARTIALMETALAREA 0.2448 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.535 2.44 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.64 -0.4 1.98 0.4 ;
      RECT 1.3 -0.4 1.64 0.575 ;
      RECT 0 -0.4 1.3 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 4.64 1.98 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
END CLKINVX3

MACRO CLKINVX2
  CLASS CORE ;
  FOREIGN CLKINVX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.98 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8124 ;
  ANTENNAPARTIALMETALAREA 0.7519 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2648 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 1.2 1.55 3.305 ;
      RECT 1.155 1.2 1.32 1.54 ;
      RECT 0.74 2.94 1.32 3.305 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4392 ;
  ANTENNAPARTIALMETALAREA 0.5575 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.6271 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 1.085 2.41 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.725 -0.4 1.98 0.4 ;
      RECT 0.385 -0.4 0.725 1.54 ;
      RECT 0 -0.4 0.385 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.45 4.64 1.98 5.44 ;
      RECT 1.07 4.395 1.45 5.44 ;
      RECT 0 4.64 1.07 5.44 ;
     END
  END VDD
END CLKINVX2

MACRO CLKINVX20
  CLASS CORE ;
  FOREIGN CLKINVX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 19.14 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 11.8547 ;
  ANTENNAPARTIALMETALAREA 16.8888 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 24.5867 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.265 2.925 18.89 3.735 ;
      RECT 16.715 1.2 18.265 3.78 ;
      RECT 15.115 1.2 16.715 1.88 ;
      RECT 16.055 2.99 16.715 3.67 ;
      RECT 15.49 2.925 16.055 3.735 ;
      RECT 14.735 2.99 15.49 3.67 ;
      RECT 13.64 1.195 15.115 1.88 ;
      RECT 14.12 2.925 14.735 3.735 ;
      RECT 13.055 2.99 14.12 3.67 ;
      RECT 10.66 1.2 13.64 1.88 ;
      RECT 12.715 2.925 13.055 3.735 ;
      RECT 11.62 2.99 12.715 3.67 ;
      RECT 11.005 2.925 11.62 3.735 ;
      RECT 10.2 2.99 11.005 3.67 ;
      RECT 10.32 1.195 10.66 1.88 ;
      RECT 8.9 1.195 10.32 1.875 ;
      RECT 9.685 2.925 10.2 3.735 ;
      RECT 8.795 2.99 9.685 3.67 ;
      RECT 8.365 2.925 8.795 3.735 ;
      RECT 7.475 2.99 8.365 3.67 ;
      RECT 7.01 2.925 7.475 3.735 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8529 ;
  ANTENNAPARTIALMETALAREA 0.2603 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.715 2.1 1.18 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.78 -0.4 19.14 0.4 ;
      RECT 15.44 -0.4 15.78 0.96 ;
      RECT 14.395 -0.4 15.44 0.4 ;
      RECT 14.055 -0.4 14.395 0.96 ;
      RECT 12.975 -0.4 14.055 0.4 ;
      RECT 12.635 -0.4 12.975 0.96 ;
      RECT 11.545 -0.4 12.635 0.4 ;
      RECT 11.205 -0.4 11.545 0.96 ;
      RECT 10.125 -0.4 11.205 0.4 ;
      RECT 9.785 -0.4 10.125 0.96 ;
      RECT 8.705 -0.4 9.785 0.4 ;
      RECT 8.365 -0.4 8.705 0.96 ;
      RECT 5.185 -0.4 8.365 0.4 ;
      RECT 4.845 -0.4 5.185 0.945 ;
      RECT 3.64 -0.4 4.845 0.4 ;
      RECT 3.3 -0.4 3.64 0.945 ;
      RECT 2.215 -0.4 3.3 0.4 ;
      RECT 1.875 -0.4 2.215 1 ;
      RECT 0 -0.4 1.875 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.015 4.64 19.14 5.44 ;
      RECT 17.675 4.12 18.015 5.44 ;
      RECT 16.59 4.64 17.675 5.44 ;
      RECT 16.25 4.12 16.59 5.44 ;
      RECT 15.17 4.64 16.25 5.44 ;
      RECT 14.83 4.12 15.17 5.44 ;
      RECT 13.745 4.64 14.83 5.44 ;
      RECT 13.405 4.12 13.745 5.44 ;
      RECT 12.335 4.64 13.405 5.44 ;
      RECT 11.995 4.12 12.335 5.44 ;
      RECT 10.915 4.64 11.995 5.44 ;
      RECT 10.575 4.065 10.915 5.44 ;
      RECT 9.48 4.64 10.575 5.44 ;
      RECT 9.14 4.065 9.48 5.44 ;
      RECT 8.06 4.64 9.14 5.44 ;
      RECT 7.72 4.065 8.06 5.44 ;
      RECT 6.64 4.64 7.72 5.44 ;
      RECT 6.3 4.075 6.64 5.44 ;
      RECT 5.07 4.64 6.3 5.44 ;
      RECT 4.73 4.06 5.07 5.44 ;
      RECT 3.635 4.64 4.73 5.44 ;
      RECT 3.295 4.06 3.635 5.44 ;
      RECT 2.165 4.64 3.295 5.44 ;
      RECT 1.825 4.09 2.165 5.44 ;
      RECT 0.805 4.64 1.825 5.44 ;
      RECT 0.465 3.05 0.805 5.44 ;
      RECT 0 4.64 0.465 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.345 2.12 16.205 2.69 ;
      RECT 5.805 1.18 6.345 3.45 ;
      RECT 5.7 1.18 5.805 3.675 ;
      RECT 2.59 1.18 5.7 1.825 ;
      RECT 5.465 2.805 5.7 3.675 ;
      RECT 4.345 2.805 5.465 3.45 ;
      RECT 2.365 2.1 5.055 2.44 ;
      RECT 4.005 2.805 4.345 3.735 ;
      RECT 2.925 2.805 4.005 3.45 ;
      RECT 2.59 2.805 2.925 3.735 ;
      RECT 2.585 2.925 2.59 3.735 ;
      RECT 1.64 2.155 2.365 2.385 ;
      RECT 1.41 1.44 1.64 3.315 ;
      RECT 1.225 1.44 1.41 1.78 ;
      RECT 1.235 2.975 1.41 3.315 ;
  END
END CLKINVX20

MACRO CLKINVX1
  CLASS CORE ;
  FOREIGN CLKINVX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.98 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.84 ;
  ANTENNAPARTIALMETALAREA 1.1746 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5245 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.485 1.82 1.83 3.22 ;
      RECT 1.255 1.35 1.485 3.885 ;
      RECT 1.04 1.35 1.255 1.855 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.316 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.19 2.38 0.925 2.81 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 -0.4 1.98 0.4 ;
      RECT 0.98 -0.4 1.32 0.575 ;
      RECT 0 -0.4 0.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.89 4.64 1.98 5.44 ;
      RECT 0.525 4.395 0.89 5.44 ;
      RECT 0 4.64 0.525 5.44 ;
     END
  END VDD
END CLKINVX1

MACRO CLKINVX16
  CLASS CORE ;
  FOREIGN CLKINVX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 16.5 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 9.3765 ;
  ANTENNAPARTIALMETALAREA 14.3603 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 20.6753 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.735 1.2 16.285 3.84 ;
      RECT 12.99 1.2 14.735 1.88 ;
      RECT 14.195 2.99 14.735 3.67 ;
      RECT 13.645 2.925 14.195 3.735 ;
      RECT 12.79 2.99 13.645 3.67 ;
      RECT 11.705 1.195 12.99 1.88 ;
      RECT 12.325 2.925 12.79 3.735 ;
      RECT 11.435 2.99 12.325 3.67 ;
      RECT 8.195 1.2 11.705 1.88 ;
      RECT 11.005 2.925 11.435 3.735 ;
      RECT 10.115 2.99 11.005 3.67 ;
      RECT 9.595 2.925 10.115 3.735 ;
      RECT 8.795 2.99 9.595 3.67 ;
      RECT 8.165 2.925 8.795 3.735 ;
      RECT 7.085 2.99 8.165 3.67 ;
      RECT 6.745 2.925 7.085 3.735 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.681 ;
  ANTENNAPARTIALMETALAREA 0.2603 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.715 2.1 1.18 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.655 -0.4 16.5 0.4 ;
      RECT 13.315 -0.4 13.655 0.96 ;
      RECT 12.27 -0.4 13.315 0.4 ;
      RECT 11.93 -0.4 12.27 0.96 ;
      RECT 10.85 -0.4 11.93 0.4 ;
      RECT 10.51 -0.4 10.85 0.96 ;
      RECT 9.42 -0.4 10.51 0.4 ;
      RECT 9.08 -0.4 9.42 0.96 ;
      RECT 8 -0.4 9.08 0.4 ;
      RECT 7.66 -0.4 8 0.96 ;
      RECT 3.64 -0.4 7.66 0.4 ;
      RECT 3.3 -0.4 3.64 1.02 ;
      RECT 2.215 -0.4 3.3 0.4 ;
      RECT 1.875 -0.4 2.215 1 ;
      RECT 0 -0.4 1.875 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.24 4.64 16.5 5.44 ;
      RECT 15.9 4.12 16.24 5.44 ;
      RECT 14.905 4.64 15.9 5.44 ;
      RECT 14.565 4.12 14.905 5.44 ;
      RECT 13.48 4.64 14.565 5.44 ;
      RECT 13.14 4.12 13.48 5.44 ;
      RECT 12.07 4.64 13.14 5.44 ;
      RECT 11.73 4.12 12.07 5.44 ;
      RECT 10.65 4.64 11.73 5.44 ;
      RECT 10.31 4.065 10.65 5.44 ;
      RECT 9.215 4.64 10.31 5.44 ;
      RECT 8.875 4.065 9.215 5.44 ;
      RECT 7.795 4.64 8.875 5.44 ;
      RECT 7.455 4.065 7.795 5.44 ;
      RECT 6.375 4.64 7.455 5.44 ;
      RECT 6.035 4.075 6.375 5.44 ;
      RECT 5.07 4.64 6.035 5.44 ;
      RECT 4.73 4.06 5.07 5.44 ;
      RECT 3.635 4.64 4.73 5.44 ;
      RECT 3.295 4.06 3.635 5.44 ;
      RECT 2.165 4.64 3.295 5.44 ;
      RECT 1.825 4.09 2.165 5.44 ;
      RECT 0.805 4.64 1.825 5.44 ;
      RECT 0.465 3.05 0.805 5.44 ;
      RECT 0 4.64 0.465 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.44 2.19 14.3 2.53 ;
      RECT 6.02 2.21 6.44 2.51 ;
      RECT 5.34 1.34 6.02 3.39 ;
      RECT 2.585 1.34 5.34 1.87 ;
      RECT 4.345 2.7 5.34 3.39 ;
      RECT 2.275 2.1 4.965 2.44 ;
      RECT 4.005 2.7 4.345 3.735 ;
      RECT 2.925 2.7 4.005 3.39 ;
      RECT 2.585 2.7 2.925 3.735 ;
      RECT 1.64 2.155 2.275 2.385 ;
      RECT 1.41 1.44 1.64 3.315 ;
      RECT 1.225 1.44 1.41 1.78 ;
      RECT 1.235 2.975 1.41 3.315 ;
  END
END CLKINVX16

MACRO CLKINVX12
  CLASS CORE ;
  FOREIGN CLKINVX12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.54 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKINVXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 6.9791 ;
  ANTENNAPARTIALMETALAREA 10.4289 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 14.5644 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.775 1.195 12.325 3.78 ;
      RECT 7.02 1.195 10.775 1.875 ;
      RECT 10.115 2.99 10.775 3.67 ;
      RECT 9.685 2.925 10.115 3.735 ;
      RECT 8.795 2.99 9.685 3.67 ;
      RECT 8.295 2.925 8.795 3.735 ;
      RECT 7.475 2.99 8.295 3.67 ;
      RECT 6.865 2.925 7.475 3.735 ;
      RECT 5.785 2.99 6.865 3.67 ;
      RECT 5.445 2.925 5.785 3.735 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5166 ;
  ANTENNAPARTIALMETALAREA 0.3331 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2243 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.51 2.1 1.105 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.925 -0.4 12.54 0.4 ;
      RECT 10.585 -0.4 10.925 0.96 ;
      RECT 9.495 -0.4 10.585 0.4 ;
      RECT 9.155 -0.4 9.495 0.96 ;
      RECT 8.075 -0.4 9.155 0.4 ;
      RECT 7.735 -0.4 8.075 0.96 ;
      RECT 6.68 -0.4 7.735 0.4 ;
      RECT 6.34 -0.4 6.68 0.96 ;
      RECT 3.55 -0.4 6.34 0.4 ;
      RECT 3.21 -0.4 3.55 1.02 ;
      RECT 0.695 -0.4 3.21 0.4 ;
      RECT 0.355 -0.4 0.695 1.685 ;
      RECT 0 -0.4 0.355 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.2 4.64 12.54 5.44 ;
      RECT 11.86 4.12 12.2 5.44 ;
      RECT 10.765 4.64 11.86 5.44 ;
      RECT 10.425 4.12 10.765 5.44 ;
      RECT 9.35 4.64 10.425 5.44 ;
      RECT 9.01 4.065 9.35 5.44 ;
      RECT 7.915 4.64 9.01 5.44 ;
      RECT 7.575 4.065 7.915 5.44 ;
      RECT 6.495 4.64 7.575 5.44 ;
      RECT 6.155 4.065 6.495 5.44 ;
      RECT 5.09 4.64 6.155 5.44 ;
      RECT 4.75 4.075 5.09 5.44 ;
      RECT 3.545 4.64 4.75 5.44 ;
      RECT 3.205 4.06 3.545 5.44 ;
      RECT 2.075 4.64 3.205 5.44 ;
      RECT 1.735 4.09 2.075 5.44 ;
      RECT 0.675 4.64 1.735 5.44 ;
      RECT 0.335 2.89 0.675 5.44 ;
      RECT 0 4.64 0.335 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.1 2.19 10.41 2.53 ;
      RECT 4.8 1.42 5.1 3.245 ;
      RECT 4.25 1.42 4.8 1.72 ;
      RECT 4.255 2.945 4.8 3.245 ;
      RECT 2.06 2.1 4.28 2.44 ;
      RECT 3.915 2.925 4.255 3.735 ;
      RECT 2.5 1.42 4.25 1.76 ;
      RECT 2.835 2.925 3.915 3.265 ;
      RECT 2.495 2.925 2.835 3.735 ;
      RECT 1.64 2.155 2.06 2.385 ;
      RECT 1.485 1.305 1.64 3.26 ;
      RECT 1.415 1.305 1.485 3.315 ;
      RECT 1.41 1.25 1.415 3.315 ;
      RECT 1.075 1.25 1.41 1.59 ;
      RECT 1.145 2.975 1.41 3.315 ;
  END
END CLKINVX12

MACRO CLKBUFXL
  CLASS CORE ;
  FOREIGN CLKBUFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6864 ;
  ANTENNAPARTIALMETALAREA 0.7833 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6994 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.195 1.22 2.425 2.99 ;
      RECT 1.92 1.22 2.195 1.45 ;
      RECT 2.12 2.635 2.195 2.99 ;
      RECT 1.88 2.76 2.12 2.99 ;
      RECT 1.58 1.11 1.92 1.45 ;
      RECT 1.54 2.76 1.88 3.1 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.108 ;
  ANTENNAPARTIALMETALAREA 0.3283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.81 2.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.12 -0.4 2.64 0.4 ;
      RECT 0.78 -0.4 1.12 0.575 ;
      RECT 0 -0.4 0.78 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.22 4.64 2.64 5.44 ;
      RECT 0.88 4.465 1.22 5.44 ;
      RECT 0 4.64 0.88 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.27 1.82 1.52 2.16 ;
      RECT 1.04 1.22 1.27 2.99 ;
      RECT 0.52 1.22 1.04 1.45 ;
      RECT 0.52 2.76 1.04 2.99 ;
      RECT 0.18 1.11 0.52 1.45 ;
      RECT 0.18 2.76 0.52 3.1 ;
  END
END CLKBUFXL

MACRO CLKBUFX8
  CLASS CORE ;
  FOREIGN CLKBUFX8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.321 ;
  ANTENNAPARTIALMETALAREA 3.168 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9714 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4 1.82 4.405 3.22 ;
      RECT 2.855 1.35 4 3.22 ;
      RECT 2.78 1.35 2.855 1.85 ;
      RECT 2.78 2.625 2.855 3.18 ;
      RECT 2.26 1.35 2.78 1.69 ;
      RECT 2.18 2.84 2.78 3.18 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6114 ;
  ANTENNAPARTIALMETALAREA 0.3121 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3833 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 1.99 1.39 2.33 ;
      RECT 0.875 1.845 1.105 2.33 ;
      RECT 0.57 1.99 0.875 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.24 -0.4 4.62 0.4 ;
      RECT 2.9 -0.4 3.24 0.965 ;
      RECT 1.96 -0.4 2.9 0.4 ;
      RECT 1.62 -0.4 1.96 0.965 ;
      RECT 0 -0.4 1.62 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.44 4.64 4.62 5.44 ;
      RECT 4.1 3.62 4.44 5.44 ;
      RECT 3.16 4.64 4.1 5.44 ;
      RECT 2.82 3.62 3.16 5.44 ;
      RECT 1.84 4.64 2.82 5.44 ;
      RECT 1.5 4.465 1.84 5.44 ;
      RECT 0.52 4.64 1.5 5.44 ;
      RECT 0.18 3.48 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.95 2.18 2.55 2.52 ;
      RECT 1.72 1.26 1.95 2.99 ;
      RECT 1.24 1.26 1.72 1.49 ;
      RECT 1.16 2.76 1.72 2.99 ;
      RECT 0.9 1.15 1.24 1.49 ;
      RECT 0.82 2.76 1.16 3.1 ;
  END
END CLKBUFX8

MACRO CLKBUFX4
  CLASS CORE ;
  FOREIGN CLKBUFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3176 ;
  ANTENNAPARTIALMETALAREA 0.887 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2542 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.35 1.26 2.5 2.66 ;
      RECT 2.12 1.26 2.35 3 ;
      RECT 1.7 1.39 2.12 1.73 ;
      RECT 2.04 2.77 2.12 3 ;
      RECT 1.7 2.77 2.04 3.11 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.288 ;
  ANTENNAPARTIALMETALAREA 0.3852 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3197 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.81 2.395 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.8 -0.4 3.3 0.4 ;
      RECT 2.46 -0.4 2.8 0.575 ;
      RECT 1.18 -0.4 2.46 0.4 ;
      RECT 0.84 -0.4 1.18 0.575 ;
      RECT 0 -0.4 0.84 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.8 4.64 3.3 5.44 ;
      RECT 2.46 4.465 2.8 5.44 ;
      RECT 1.28 4.64 2.46 5.44 ;
      RECT 1.225 4.465 1.28 5.44 ;
      RECT 0.995 4.41 1.225 5.44 ;
      RECT 0.94 4.465 0.995 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.27 2.06 1.89 2.4 ;
      RECT 1.04 1.36 1.27 2.97 ;
      RECT 0.52 1.36 1.04 1.59 ;
      RECT 0.52 2.74 1.04 2.97 ;
      RECT 0.18 1.25 0.52 1.59 ;
      RECT 0.18 2.74 0.52 3.08 ;
  END
END CLKBUFX4

MACRO CLKBUFX3
  CLASS CORE ;
  FOREIGN CLKBUFX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.9927 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5917 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.77 1.205 1.88 1.545 ;
      RECT 1.77 1.82 1.84 3.16 ;
      RECT 1.54 1.205 1.77 3.16 ;
      RECT 1.5 1.82 1.54 3.16 ;
      RECT 1.46 1.82 1.5 2.66 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2232 ;
  ANTENNAPARTIALMETALAREA 0.2241 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0123 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.555 2.36 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.46 -0.4 2.64 0.4 ;
      RECT 2.12 -0.4 2.46 0.575 ;
      RECT 1.18 -0.4 2.12 0.4 ;
      RECT 0.84 -0.4 1.18 0.575 ;
      RECT 0 -0.4 0.84 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.46 4.64 2.64 5.44 ;
      RECT 2.12 4.465 2.46 5.44 ;
      RECT 1.195 4.64 2.12 5.44 ;
      RECT 0.81 4.465 1.195 5.44 ;
      RECT 0 4.64 0.81 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.115 1.975 1.225 2.315 ;
      RECT 0.885 1.135 1.115 3.155 ;
      RECT 0.52 1.135 0.885 1.365 ;
      RECT 0.52 2.925 0.885 3.155 ;
      RECT 0.18 1.025 0.52 1.365 ;
      RECT 0.18 2.925 0.52 3.265 ;
  END
END CLKBUFX3

MACRO CLKBUFX2
  CLASS CORE ;
  FOREIGN CLKBUFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2 ;
  ANTENNAPARTIALMETALAREA 0.7946 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5139 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.2 1.265 2.425 2.98 ;
      RECT 2.195 1.155 2.2 2.98 ;
      RECT 1.64 1.155 2.195 1.495 ;
      RECT 2.12 2.635 2.195 3.09 ;
      RECT 1.6 2.75 2.12 3.09 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1944 ;
  ANTENNAPARTIALMETALAREA 0.3838 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3409 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.9 2.26 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.22 -0.4 2.64 0.4 ;
      RECT 0.88 -0.4 1.22 0.575 ;
      RECT 0 -0.4 0.88 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 1.125 4.465 1.18 5.44 ;
      RECT 0.895 4.41 1.125 5.44 ;
      RECT 0.84 4.465 0.895 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.37 2.06 1.62 2.4 ;
      RECT 1.14 1.265 1.37 2.98 ;
      RECT 0.62 1.265 1.14 1.495 ;
      RECT 0.62 2.75 1.14 2.98 ;
      RECT 0.28 1.155 0.62 1.495 ;
      RECT 0.28 2.75 0.62 3.09 ;
  END
END CLKBUFX2

MACRO CLKBUFX20
  CLASS CORE ;
  FOREIGN CLKBUFX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 8.8679 ;
  ANTENNAPARTIALMETALAREA 18.1738 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 23.0391 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.76 1.2 14.965 3.84 ;
      RECT 13.415 1.125 14.76 3.84 ;
      RECT 4.7 1.125 13.415 1.925 ;
      RECT 13.34 2.66 13.415 3.525 ;
      RECT 4.66 2.725 13.34 3.525 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.5326 ;
  ANTENNAPARTIALMETALAREA 1.1077 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8637 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.085 1.99 3.74 2.33 ;
      RECT 2.855 1.845 3.085 2.33 ;
      RECT 0.58 1.99 2.855 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.8 -0.4 15.84 0.4 ;
      RECT 10.46 -0.4 10.8 0.895 ;
      RECT 9.52 -0.4 10.46 0.4 ;
      RECT 9.18 -0.4 9.52 0.895 ;
      RECT 8.24 -0.4 9.18 0.4 ;
      RECT 7.9 -0.4 8.24 0.895 ;
      RECT 6.96 -0.4 7.9 0.4 ;
      RECT 6.62 -0.4 6.96 0.895 ;
      RECT 5.68 -0.4 6.62 0.4 ;
      RECT 5.34 -0.4 5.68 0.895 ;
      RECT 4.4 -0.4 5.34 0.4 ;
      RECT 4.06 -0.4 4.4 0.96 ;
      RECT 2.96 -0.4 4.06 0.4 ;
      RECT 2.62 -0.4 2.96 0.96 ;
      RECT 1.52 -0.4 2.62 0.4 ;
      RECT 1.18 -0.4 1.52 0.96 ;
      RECT 0 -0.4 1.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.64 4.64 15.84 5.44 ;
      RECT 14.585 4.465 14.64 5.44 ;
      RECT 14.355 4.41 14.585 5.44 ;
      RECT 14.3 4.465 14.355 5.44 ;
      RECT 13.32 4.64 14.3 5.44 ;
      RECT 12.98 4.09 13.32 5.44 ;
      RECT 12.04 4.64 12.98 5.44 ;
      RECT 11.7 4.09 12.04 5.44 ;
      RECT 10.76 4.64 11.7 5.44 ;
      RECT 10.42 4.09 10.76 5.44 ;
      RECT 9.48 4.64 10.42 5.44 ;
      RECT 9.14 4.09 9.48 5.44 ;
      RECT 8.2 4.64 9.14 5.44 ;
      RECT 7.86 4.09 8.2 5.44 ;
      RECT 6.92 4.64 7.86 5.44 ;
      RECT 6.58 4.02 6.92 5.44 ;
      RECT 5.64 4.64 6.58 5.44 ;
      RECT 5.3 4.02 5.64 5.44 ;
      RECT 4.36 4.64 5.3 5.44 ;
      RECT 4.02 3.945 4.36 5.44 ;
      RECT 3.08 4.64 4.02 5.44 ;
      RECT 2.74 3.945 3.08 5.44 ;
      RECT 1.8 4.64 2.74 5.44 ;
      RECT 1.46 3.945 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.945 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.42 2.155 12.92 2.495 ;
      RECT 4.08 1.19 4.42 3.18 ;
      RECT 1.9 1.19 4.08 1.53 ;
      RECT 0.82 2.84 4.08 3.18 ;
  END
END CLKBUFX20

MACRO CLKBUFX1
  CLASS CORE ;
  FOREIGN CLKBUFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6964 ;
  ANTENNAPARTIALMETALAREA 0.8108 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8054 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.195 1.22 2.425 3.05 ;
      RECT 1.92 1.22 2.195 1.45 ;
      RECT 2.12 2.635 2.195 3.05 ;
      RECT 1.84 2.82 2.12 3.05 ;
      RECT 1.58 1.11 1.92 1.45 ;
      RECT 1.5 2.82 1.84 3.16 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2304 ;
  ANTENNAPARTIALMETALAREA 0.3283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.81 2.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.12 -0.4 2.64 0.4 ;
      RECT 0.78 -0.4 1.12 0.575 ;
      RECT 0 -0.4 0.78 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 0.84 4.465 1.18 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.27 2.06 1.52 2.4 ;
      RECT 1.04 1.22 1.27 2.99 ;
      RECT 0.52 1.22 1.04 1.45 ;
      RECT 0.52 2.76 1.04 2.99 ;
      RECT 0.18 1.11 0.52 1.45 ;
      RECT 0.18 2.76 0.52 3.1 ;
  END
END CLKBUFX1

MACRO CLKBUFX16
  CLASS CORE ;
  FOREIGN CLKBUFX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.54 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 7.7705 ;
  ANTENNAPARTIALMETALAREA 14.8938 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 18.6931 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.12 1.2 12.325 3.84 ;
      RECT 10.775 1.125 12.12 3.84 ;
      RECT 4.06 1.125 10.775 1.925 ;
      RECT 10.7 2.66 10.775 3.525 ;
      RECT 4.12 2.725 10.7 3.525 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.8312 ;
  ANTENNAPARTIALMETALAREA 0.595 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2154 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.28 1.79 3.03 2.13 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.08 -0.4 12.54 0.4 ;
      RECT 8.74 -0.4 9.08 0.895 ;
      RECT 7.64 -0.4 8.74 0.4 ;
      RECT 7.3 -0.4 7.64 0.895 ;
      RECT 6.32 -0.4 7.3 0.4 ;
      RECT 5.98 -0.4 6.32 0.895 ;
      RECT 5.04 -0.4 5.98 0.4 ;
      RECT 4.7 -0.4 5.04 0.895 ;
      RECT 3.76 -0.4 4.7 0.4 ;
      RECT 3.42 -0.4 3.76 0.895 ;
      RECT 2.32 -0.4 3.42 0.4 ;
      RECT 1.98 -0.4 2.32 0.895 ;
      RECT 0 -0.4 1.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.58 4.64 12.54 5.44 ;
      RECT 11.24 4.09 11.58 5.44 ;
      RECT 10.26 4.64 11.24 5.44 ;
      RECT 9.92 4.02 10.26 5.44 ;
      RECT 8.98 4.64 9.92 5.44 ;
      RECT 8.64 4.02 8.98 5.44 ;
      RECT 7.7 4.64 8.64 5.44 ;
      RECT 7.36 4.02 7.7 5.44 ;
      RECT 6.38 4.64 7.36 5.44 ;
      RECT 6.04 4.02 6.38 5.44 ;
      RECT 5.1 4.64 6.04 5.44 ;
      RECT 4.76 4.02 5.1 5.44 ;
      RECT 3.82 4.64 4.76 5.44 ;
      RECT 3.48 4.02 3.82 5.44 ;
      RECT 2.5 4.64 3.48 5.44 ;
      RECT 2.16 3.62 2.5 5.44 ;
      RECT 1.18 4.64 2.16 5.44 ;
      RECT 1.125 4.465 1.18 5.44 ;
      RECT 0.895 4.41 1.125 5.44 ;
      RECT 0.84 4.465 0.895 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.78 2.155 10.36 2.495 ;
      RECT 3.44 1.15 3.78 3.1 ;
      RECT 1.26 1.15 3.44 1.49 ;
      RECT 1.52 2.76 3.44 3.1 ;
  END
END CLKBUFX16

MACRO CLKBUFX12
  CLASS CORE ;
  FOREIGN CLKBUFX12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CLKBUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 5.484 ;
  ANTENNAPARTIALMETALAREA 9.7582 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 13.939 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.48 1.2 9.685 3.28 ;
      RECT 8.135 1.18 9.48 3.35 ;
      RECT 3.46 1.18 8.135 1.86 ;
      RECT 8.06 2.66 8.135 3.35 ;
      RECT 3.38 2.67 8.06 3.35 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.5372 ;
  ANTENNAPARTIALMETALAREA 0.7065 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6129 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.99 2.58 2.33 ;
      RECT 1.535 1.845 1.765 2.33 ;
      RECT 0.6 1.99 1.535 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7 -0.4 10.56 0.4 ;
      RECT 6.66 -0.4 7 0.95 ;
      RECT 5.72 -0.4 6.66 0.4 ;
      RECT 5.38 -0.4 5.72 0.95 ;
      RECT 4.44 -0.4 5.38 0.4 ;
      RECT 4.1 -0.4 4.44 0.95 ;
      RECT 3.16 -0.4 4.1 0.4 ;
      RECT 2.82 -0.4 3.16 0.95 ;
      RECT 1.88 -0.4 2.82 0.4 ;
      RECT 1.54 -0.4 1.88 0.95 ;
      RECT 0 -0.4 1.54 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.52 4.64 10.56 5.44 ;
      RECT 9.465 4.465 9.52 5.44 ;
      RECT 9.235 4.41 9.465 5.44 ;
      RECT 9.18 4.465 9.235 5.44 ;
      RECT 8.2 4.64 9.18 5.44 ;
      RECT 7.86 3.675 8.2 5.44 ;
      RECT 6.92 4.64 7.86 5.44 ;
      RECT 6.58 3.675 6.92 5.44 ;
      RECT 5.64 4.64 6.58 5.44 ;
      RECT 5.3 3.675 5.64 5.44 ;
      RECT 4.36 4.64 5.3 5.44 ;
      RECT 4.02 3.675 4.36 5.44 ;
      RECT 3.08 4.64 4.02 5.44 ;
      RECT 2.74 3.725 3.08 5.44 ;
      RECT 1.8 4.64 2.74 5.44 ;
      RECT 1.46 3.705 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.705 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.15 2.09 7.8 2.43 ;
      RECT 2.81 1.34 3.15 3.1 ;
      RECT 2.18 1.34 2.81 1.68 ;
      RECT 0.82 2.76 2.81 3.1 ;
  END
END CLKBUFX12

MACRO BUFXL
  CLASS CORE ;
  FOREIGN BUFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5216 ;
  ANTENNAPARTIALMETALAREA 0.8361 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.195 1.15 2.425 3.05 ;
      RECT 1.88 1.15 2.195 1.38 ;
      RECT 2.12 2.635 2.195 3.05 ;
      RECT 1.84 2.82 2.12 3.05 ;
      RECT 1.54 1.04 1.88 1.38 ;
      RECT 1.5 2.82 1.84 3.16 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.81 2.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.12 -0.4 2.64 0.4 ;
      RECT 0.78 -0.4 1.12 0.575 ;
      RECT 0 -0.4 0.78 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 0.84 4.465 1.18 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.27 2.06 1.52 2.4 ;
      RECT 1.04 1.22 1.27 2.99 ;
      RECT 0.52 1.22 1.04 1.45 ;
      RECT 0.52 2.76 1.04 2.99 ;
      RECT 0.18 1.11 0.52 1.45 ;
      RECT 0.18 2.76 0.52 3.1 ;
  END
END BUFXL

MACRO NBUFFX8_LVT
  CLASS CORE ;
  FOREIGN NBUFFX8_LVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.6056 ;
  ANTENNAPARTIALMETALAREA 3.8231 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.466 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.53 1.82 5.065 3.22 ;
      RECT 4.2 1.82 4.53 3.25 ;
      RECT 3.515 1.29 4.2 3.25 ;
      RECT 3.44 1.29 3.515 1.85 ;
      RECT 3.44 2.63 3.515 3.25 ;
      RECT 2.26 1.29 3.44 1.77 ;
      RECT 2.18 2.77 3.44 3.25 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8634 ;
  ANTENNAPARTIALMETALAREA 0.3087 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3727 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 1.99 1.38 2.33 ;
      RECT 0.875 1.845 1.105 2.33 ;
      RECT 0.57 1.99 0.875 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.52 -0.4 5.94 0.4 ;
      RECT 4.18 -0.4 4.52 0.95 ;
      RECT 3.24 -0.4 4.18 0.4 ;
      RECT 2.9 -0.4 3.24 0.95 ;
      RECT 1.96 -0.4 2.9 0.4 ;
      RECT 1.62 -0.4 1.96 0.895 ;
      RECT 0.52 -0.4 1.62 0.4 ;
      RECT 0.18 -0.4 0.52 0.95 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.44 4.64 5.94 5.44 ;
      RECT 4.1 3.62 4.44 5.44 ;
      RECT 3.16 4.64 4.1 5.44 ;
      RECT 2.82 3.62 3.16 5.44 ;
      RECT 1.88 4.64 2.82 5.44 ;
      RECT 1.54 3.705 1.88 5.44 ;
      RECT 0.6 4.64 1.54 5.44 ;
      RECT 0.26 3.705 0.6 5.44 ;
      RECT 0 4.64 0.26 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.95 2.18 3.21 2.52 ;
      RECT 1.61 1.15 1.95 3.1 ;
      RECT 0.9 1.15 1.61 1.49 ;
      RECT 0.9 2.76 1.61 3.1 ;
  END
END NBUFFX8_LVT

MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5984 ;
  ANTENNAPARTIALMETALAREA 1.4894 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5792 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.2 1.26 2.5 3.08 ;
      RECT 2.12 1.26 2.2 3.22 ;
      RECT 2.04 1.26 2.12 1.73 ;
      RECT 2.04 2.74 2.12 3.22 ;
      RECT 1.7 0.92 2.04 1.73 ;
      RECT 1.7 2.74 2.04 4.02 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.432 ;
  ANTENNAPARTIALMETALAREA 0.3795 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.8 2.395 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.8 -0.4 3.3 0.4 ;
      RECT 2.46 -0.4 2.8 0.575 ;
      RECT 1.28 -0.4 2.46 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.8 4.64 3.3 5.44 ;
      RECT 2.46 3.94 2.8 5.44 ;
      RECT 1.28 4.64 2.46 5.44 ;
      RECT 0.94 3.94 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.38 2.005 1.89 2.455 ;
      RECT 1.04 1.25 1.38 3.08 ;
      RECT 0.52 1.25 1.04 1.59 ;
      RECT 0.52 2.74 1.04 3.08 ;
      RECT 0.18 0.78 0.52 1.59 ;
      RECT 0.18 2.74 0.52 4.02 ;
  END
END BUFX4

MACRO BUFX3
  CLASS CORE ;
  FOREIGN BUFX3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2324 ;
  ANTENNAPARTIALMETALAREA 0.668 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5917 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.77 1.205 1.88 1.545 ;
      RECT 1.77 1.82 1.84 3.16 ;
      RECT 1.54 1.205 1.77 3.16 ;
      RECT 1.5 1.82 1.54 3.16 ;
      RECT 1.46 1.82 1.5 2.66 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.324 ;
  ANTENNAPARTIALMETALAREA 0.224 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0123 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.555 2.36 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.44 -0.4 2.64 0.4 ;
      RECT 2.1 -0.4 2.44 0.575 ;
      RECT 0 -0.4 2.1 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.08 4.64 2.64 5.44 ;
      RECT 0.74 4.465 1.08 5.44 ;
      RECT 0 4.64 0.74 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.115 1.975 1.225 2.315 ;
      RECT 0.885 1.135 1.115 3.155 ;
      RECT 0.52 1.135 0.885 1.365 ;
      RECT 0.52 2.925 0.885 3.155 ;
      RECT 0.18 1.025 0.52 1.365 ;
      RECT 0.18 2.925 0.52 3.265 ;
  END
END BUFX3

MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.48 ;
  ANTENNAPARTIALMETALAREA 0.6624 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1853 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.35 1.845 2.425 2.075 ;
      RECT 2.12 1.5 2.35 2.98 ;
      RECT 1.98 1.5 2.12 1.73 ;
      RECT 1.94 2.75 2.12 2.98 ;
      RECT 1.64 1.39 1.98 1.73 ;
      RECT 1.6 2.75 1.94 3.09 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.216 ;
  ANTENNAPARTIALMETALAREA 0.3787 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3303 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.89 2.26 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.22 -0.4 2.64 0.4 ;
      RECT 0.88 -0.4 1.22 0.575 ;
      RECT 0 -0.4 0.88 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 1.125 4.465 1.18 5.44 ;
      RECT 0.895 4.41 1.125 5.44 ;
      RECT 0.84 4.465 0.895 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.37 2.06 1.62 2.4 ;
      RECT 1.14 1.265 1.37 2.99 ;
      RECT 0.62 1.265 1.14 1.495 ;
      RECT 0.62 2.76 1.14 2.99 ;
      RECT 0.28 1.155 0.62 1.495 ;
      RECT 0.28 2.76 0.62 3.1 ;
  END
END BUFX2

MACRO BUFX20
  CLASS CORE ;
  FOREIGN BUFX20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.56 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 6.5045 ;
  ANTENNAPARTIALMETALAREA 12.8451 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 15.9583 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.795 1.125 10.345 3.84 ;
      RECT 3.42 1.125 8.795 1.925 ;
      RECT 8.72 2.66 8.795 3.525 ;
      RECT 3.38 2.725 8.72 3.525 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.1792 ;
  ANTENNAPARTIALMETALAREA 0.6283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.3691 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.99 2.5 2.33 ;
      RECT 1.535 1.845 1.765 2.33 ;
      RECT 0.75 1.99 1.535 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.56 -0.4 10.56 0.4 ;
      RECT 9.22 -0.4 9.56 0.575 ;
      RECT 8.24 -0.4 9.22 0.4 ;
      RECT 7.9 -0.4 8.24 0.895 ;
      RECT 6.96 -0.4 7.9 0.4 ;
      RECT 6.62 -0.4 6.96 0.895 ;
      RECT 5.68 -0.4 6.62 0.4 ;
      RECT 5.34 -0.4 5.68 0.895 ;
      RECT 4.4 -0.4 5.34 0.4 ;
      RECT 4.06 -0.4 4.4 0.895 ;
      RECT 3.12 -0.4 4.06 0.4 ;
      RECT 2.78 -0.4 3.12 0.965 ;
      RECT 1.8 -0.4 2.78 0.4 ;
      RECT 1.46 -0.4 1.8 1.045 ;
      RECT 0.52 -0.4 1.46 0.4 ;
      RECT 0.18 -0.4 0.52 1.045 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 9.52 4.64 10.56 5.44 ;
      RECT 9.465 4.465 9.52 5.44 ;
      RECT 9.235 4.41 9.465 5.44 ;
      RECT 9.18 4.465 9.235 5.44 ;
      RECT 8.2 4.64 9.18 5.44 ;
      RECT 7.86 4.09 8.2 5.44 ;
      RECT 6.92 4.64 7.86 5.44 ;
      RECT 6.58 4.09 6.92 5.44 ;
      RECT 5.64 4.64 6.58 5.44 ;
      RECT 5.3 4.02 5.64 5.44 ;
      RECT 4.36 4.64 5.3 5.44 ;
      RECT 4.02 4.02 4.36 5.44 ;
      RECT 3.08 4.64 4.02 5.44 ;
      RECT 2.74 3.605 3.08 5.44 ;
      RECT 1.8 4.64 2.74 5.44 ;
      RECT 1.46 3.605 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.605 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.145 2.155 8.26 2.495 ;
      RECT 2.805 1.345 3.145 3.18 ;
      RECT 2.1 1.345 2.805 1.685 ;
      RECT 0.82 2.84 2.805 3.18 ;
      RECT 1.16 1.345 2.1 1.575 ;
      RECT 0.82 1.345 1.16 1.685 ;
  END
END BUFX20

MACRO BUFX1
  CLASS CORE ;
  FOREIGN BUFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.75 ;
  ANTENNAPARTIALMETALAREA 0.8361 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.922 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.195 1.15 2.425 3.05 ;
      RECT 1.88 1.15 2.195 1.38 ;
      RECT 2.12 2.635 2.195 3.05 ;
      RECT 1.84 2.82 2.12 3.05 ;
      RECT 1.54 1.04 1.88 1.38 ;
      RECT 1.5 2.82 1.84 3.16 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.3283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.755 0.81 2.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.12 -0.4 2.64 0.4 ;
      RECT 0.78 -0.4 1.12 0.575 ;
      RECT 0 -0.4 0.78 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 0.84 4.465 1.18 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.27 2.06 1.52 2.4 ;
      RECT 1.04 1.22 1.27 2.99 ;
      RECT 0.52 1.22 1.04 1.45 ;
      RECT 0.52 2.76 1.04 2.99 ;
      RECT 0.18 1.11 0.52 1.45 ;
      RECT 0.18 2.76 0.52 3.1 ;
  END
END BUFX1

MACRO BUFX16
  CLASS CORE ;
  FOREIGN BUFX16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.58 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 5.2896 ;
  ANTENNAPARTIALMETALAREA 10.1597 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 12.3967 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.815 1.125 8.365 3.84 ;
      RECT 2.78 1.125 6.815 1.925 ;
      RECT 6.74 2.625 6.815 3.525 ;
      RECT 3.42 2.725 6.74 3.525 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.7295 ;
  ANTENNAPARTIALMETALAREA 0.5205 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0193 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 2.19 2.04 2.53 ;
      RECT 1.535 2.19 1.765 2.635 ;
      RECT 0.58 2.19 1.535 2.53 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.72 -0.4 8.58 0.4 ;
      RECT 7.38 -0.4 7.72 0.575 ;
      RECT 6.36 -0.4 7.38 0.4 ;
      RECT 6.02 -0.4 6.36 0.895 ;
      RECT 5.04 -0.4 6.02 0.4 ;
      RECT 4.7 -0.4 5.04 0.895 ;
      RECT 3.76 -0.4 4.7 0.4 ;
      RECT 3.42 -0.4 3.76 0.895 ;
      RECT 2.44 -0.4 3.42 0.4 ;
      RECT 2.1 -0.4 2.44 0.97 ;
      RECT 1.16 -0.4 2.1 0.4 ;
      RECT 0.82 -0.4 1.16 0.965 ;
      RECT 0 -0.4 0.82 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.4 4.64 8.58 5.44 ;
      RECT 8.06 4.465 8.4 5.44 ;
      RECT 7.04 4.64 8.06 5.44 ;
      RECT 6.7 4.465 7.04 5.44 ;
      RECT 5.68 4.64 6.7 5.44 ;
      RECT 5.34 4.02 5.68 5.44 ;
      RECT 4.4 4.64 5.34 5.44 ;
      RECT 4.06 4.02 4.4 5.44 ;
      RECT 3.12 4.64 4.06 5.44 ;
      RECT 2.78 4.02 3.12 5.44 ;
      RECT 1.8 4.64 2.78 5.44 ;
      RECT 1.46 3.395 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.395 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.505 2.155 6.51 2.495 ;
      RECT 2.275 1.405 2.505 3.12 ;
      RECT 0.18 1.405 2.275 1.745 ;
      RECT 2.1 2.76 2.275 3.12 ;
      RECT 1.16 2.89 2.1 3.12 ;
      RECT 0.82 2.76 1.16 3.12 ;
  END
END BUFX16

MACRO BUFX12
  CLASS CORE ;
  FOREIGN BUFX12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BUFXL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.9084 ;
  ANTENNAPARTIALMETALAREA 4.4631 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.0772 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.835 1.26 6.385 3.22 ;
      RECT 4.76 1.35 4.835 1.85 ;
      RECT 4.76 2.63 4.835 3.18 ;
      RECT 2.82 1.35 4.76 1.69 ;
      RECT 2.74 2.84 4.76 3.18 ;
     END
  END Y

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.2927 ;
  ANTENNAPARTIALMETALAREA 0.4821 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.9133 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 1.99 2.03 2.33 ;
      RECT 0.875 1.845 1.105 2.33 ;
      RECT 0.71 1.99 0.875 2.33 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.36 -0.4 6.6 0.4 ;
      RECT 6.02 -0.4 6.36 0.95 ;
      RECT 5.08 -0.4 6.02 0.4 ;
      RECT 4.74 -0.4 5.08 0.95 ;
      RECT 3.8 -0.4 4.74 0.4 ;
      RECT 3.46 -0.4 3.8 0.965 ;
      RECT 2.52 -0.4 3.46 0.4 ;
      RECT 2.18 -0.4 2.52 0.965 ;
      RECT 1.2 -0.4 2.18 0.4 ;
      RECT 0.86 -0.4 1.2 0.575 ;
      RECT 0 -0.4 0.86 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.42 4.64 6.6 5.44 ;
      RECT 6.08 4.02 6.42 5.44 ;
      RECT 5.05 4.64 6.08 5.44 ;
      RECT 4.71 4.02 5.05 5.44 ;
      RECT 3.72 4.64 4.71 5.44 ;
      RECT 3.38 4.02 3.72 5.44 ;
      RECT 2.44 4.64 3.38 5.44 ;
      RECT 2.1 3.705 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 3.705 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.51 2.18 4.375 2.52 ;
      RECT 2.28 1.45 2.51 2.99 ;
      RECT 1.88 1.45 2.28 1.68 ;
      RECT 1.8 2.76 2.28 2.99 ;
      RECT 1.54 1.34 1.88 1.68 ;
      RECT 1.46 2.76 1.8 3.1 ;
      RECT 0.52 1.34 1.54 1.57 ;
      RECT 0.52 2.76 1.46 2.99 ;
      RECT 0.29 1.34 0.52 1.635 ;
      RECT 0.18 2.76 0.52 3.1 ;
      RECT 0.18 1.405 0.29 1.635 ;
  END
END BUFX12

MACRO AOI33XL
  CLASS CORE ;
  FOREIGN AOI33XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2132 ;
  ANTENNAPARTIALMETALAREA 1.6824 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.8864 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.835 1.24 5.065 3.45 ;
      RECT 2.11 1.24 4.835 1.47 ;
      RECT 4.56 3.22 4.835 3.45 ;
      RECT 4.22 3.22 4.56 3.56 ;
      RECT 3.12 3.22 4.22 3.45 ;
      RECT 2.78 3.22 3.12 3.56 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2499 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.685 0.63 2.195 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.3136 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.29 2.685 1.41 3.025 ;
      RECT 0.755 2.685 1.29 3.195 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2271 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.58 1.7 2.09 2.125 ;
      RECT 1.535 1.845 1.58 2.075 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2433 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.05 1.715 4.48 2.215 ;
      RECT 3.98 1.715 4.05 2.12 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2682 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.02 2.265 3.745 2.635 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2889 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1395 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.17 2.405 2.71 2.94 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.33 -0.4 5.28 0.4 ;
      RECT 3.99 -0.4 4.33 0.575 ;
      RECT 0.52 -0.4 3.99 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.64 4.64 5.28 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0.52 4.64 1.3 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.46 3.695 3.84 4.025 ;
      RECT 2.4 3.795 3.46 4.025 ;
      RECT 2.115 3.64 2.4 4.025 ;
      RECT 0.74 3.64 2.115 3.98 ;
  END
END AOI33XL

MACRO AOI33X4
  CLASS CORE ;
  FOREIGN AOI33X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI33XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3188 ;
  ANTENNAPARTIALMETALAREA 1.0438 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8478 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.97 1.82 7.12 3.22 ;
      RECT 6.74 1.43 6.97 3.22 ;
      RECT 6.405 1.43 6.74 1.66 ;
      RECT 6.065 2.82 6.74 3.16 ;
      RECT 6.065 1.32 6.405 1.66 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2137 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9805 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.65 0.615 2.1 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.3437 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2455 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.355 1.425 2.905 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.245 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.75 2.16 2.1 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2358 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.055 2.105 4.48 2.66 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.28 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.975 1.82 3.82 2.15 ;
      RECT 2.97 1.92 2.975 2.15 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2731 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.585 2.405 3.16 2.88 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.045 -0.4 7.26 0.4 ;
      RECT 6.705 -0.4 7.045 0.96 ;
      RECT 5.725 -0.4 6.705 0.4 ;
      RECT 5.385 -0.4 5.725 0.9 ;
      RECT 4.28 -0.4 5.385 0.4 ;
      RECT 3.94 -0.4 4.28 0.575 ;
      RECT 0.52 -0.4 3.94 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.045 4.64 7.26 5.44 ;
      RECT 6.705 3.68 7.045 5.44 ;
      RECT 5.765 4.64 6.705 5.44 ;
      RECT 5.425 3.87 5.765 5.44 ;
      RECT 1.645 4.64 5.425 5.44 ;
      RECT 1.305 4.465 1.645 5.44 ;
      RECT 0.525 4.64 1.305 5.44 ;
      RECT 0.185 4.465 0.525 5.44 ;
      RECT 0 4.64 0.185 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.43 2.085 6.44 2.315 ;
      RECT 5.2 1.18 5.43 3.585 ;
      RECT 5.01 1.18 5.2 1.41 ;
      RECT 5.11 3.355 5.2 3.585 ;
      RECT 4.88 3.355 5.11 4.045 ;
      RECT 4.78 0.665 5.01 1.41 ;
      RECT 4.725 1.645 4.955 3.12 ;
      RECT 4.665 3.815 4.88 4.045 ;
      RECT 4.665 0.665 4.78 0.895 ;
      RECT 4.285 1.645 4.725 1.875 ;
      RECT 4.405 2.89 4.725 3.12 ;
      RECT 4.175 2.89 4.405 3.37 ;
      RECT 4.055 1.16 4.285 1.875 ;
      RECT 3.07 3.14 4.175 3.37 ;
      RECT 2.345 1.16 4.055 1.39 ;
      RECT 3.545 3.925 3.895 4.405 ;
      RECT 2.35 3.925 3.545 4.155 ;
      RECT 2.84 3.14 3.07 3.525 ;
      RECT 2.12 3.265 2.35 4.155 ;
      RECT 2.115 1.025 2.345 1.39 ;
      RECT 0.8 3.265 2.12 3.605 ;
  END
END AOI33X4

MACRO AOI33X2
  CLASS CORE ;
  FOREIGN AOI33X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.58 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI33XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.5891 ;
  ANTENNAPARTIALMETALAREA 2.8822 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 13.4408 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.135 0.805 8.365 3.305 ;
      RECT 8.06 0.805 8.135 1.285 ;
      RECT 4.745 3.075 8.135 3.305 ;
      RECT 3.53 0.805 8.06 1.035 ;
      RECT 3.3 0.805 3.53 1.48 ;
      RECT 2.02 1.25 3.3 1.48 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 1.0388 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9555 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.615 2.85 3.995 3.19 ;
      RECT 0.7 2.96 3.615 3.19 ;
      RECT 0.47 2.405 0.7 3.19 ;
      RECT 0.215 2.405 0.47 2.635 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 0.652 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2489 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.085 2.5 3.275 2.73 ;
      RECT 2.855 1.845 3.085 2.73 ;
      RECT 1.095 2.5 2.855 2.73 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 0.2157 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.78 1.845 2.155 2.27 ;
      RECT 1.535 1.845 1.78 2.075 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 1.1522 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.5544 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.6 1.265 7.83 2.02 ;
      RECT 4.47 1.265 7.6 1.495 ;
      RECT 4.24 1.265 4.47 2.325 ;
      RECT 4.175 1.845 4.24 2.075 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 0.7716 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8001 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.77 1.725 7 2.41 ;
      RECT 5.27 1.725 6.77 1.955 ;
      RECT 5.04 1.725 5.27 2.69 ;
      RECT 4.835 2.405 5.04 2.635 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.777 ;
  ANTENNAPARTIALMETALAREA 0.323 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.75 2.205 6.46 2.66 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.005 -0.4 8.58 0.4 ;
      RECT 7.665 -0.4 8.005 0.575 ;
      RECT 4.245 -0.4 7.665 0.4 ;
      RECT 3.905 -0.4 4.245 0.575 ;
      RECT 0.52 -0.4 3.905 0.4 ;
      RECT 0.18 -0.4 0.52 1.755 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.72 4.64 8.58 5.44 ;
      RECT 3.38 4.07 3.72 5.44 ;
      RECT 2.44 4.64 3.38 5.44 ;
      RECT 2.1 4.07 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 4.07 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 7.955 3.765 8.295 4.105 ;
      RECT 7.005 3.82 7.955 4.05 ;
      RECT 6.665 3.765 7.005 4.105 ;
      RECT 5.725 3.82 6.665 4.05 ;
      RECT 5.385 3.765 5.725 4.105 ;
      RECT 4.445 3.82 5.385 4.05 ;
      RECT 4.335 3.765 4.445 4.105 ;
      RECT 4.105 3.42 4.335 4.105 ;
      RECT 0.18 3.42 4.105 3.65 ;
  END
END AOI33X2

MACRO AOI33X1
  CLASS CORE ;
  FOREIGN AOI33X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI33XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.7424 ;
  ANTENNAPARTIALMETALAREA 1.8882 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.374 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.99 2.405 5.065 2.635 ;
      RECT 4.835 0.905 4.99 3.135 ;
      RECT 4.76 0.905 4.835 3.22 ;
      RECT 2.02 0.905 4.76 1.135 ;
      RECT 4.72 2.905 4.76 3.22 ;
      RECT 4.38 2.905 4.72 3.83 ;
      RECT 3.515 2.905 4.38 3.135 ;
      RECT 2.94 2.905 3.515 3.245 ;
     END
  END Y

  PIN B2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2695 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1501 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.76 0.84 2.145 ;
     END
  END B2

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2827 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1819 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.75 2.38 1.475 2.77 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.3146 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2243 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.42 1.66 2.135 2.1 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2626 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.9 1.61 4.405 2.13 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2347 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.52 2.38 3.915 2.66 ;
      RECT 3.18 2.295 3.52 2.66 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2374 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.41 2.295 2.925 2.66 ;
      RECT 2.195 2.405 2.41 2.635 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.24 -0.4 5.28 0.4 ;
      RECT 3.9 -0.4 4.24 0.575 ;
      RECT 0.52 -0.4 3.9 0.4 ;
      RECT 0.18 -0.4 0.52 1.43 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2 4.64 5.28 5.44 ;
      RECT 1.66 4.465 2 5.44 ;
      RECT 0.52 4.64 1.66 5.44 ;
      RECT 0.18 3.01 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.66 3.61 4 4.005 ;
      RECT 2.56 3.775 3.66 4.005 ;
      RECT 2.22 3.01 2.56 4.005 ;
      RECT 1.24 3.775 2.22 4.005 ;
      RECT 0.9 3.01 1.24 4.005 ;
  END
END AOI33X1

MACRO AOI32XL
  CLASS CORE ;
  FOREIGN AOI32XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.788 ;
  ANTENNAPARTIALMETALAREA 1.3345 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.3388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.33 1.845 4.405 2.075 ;
      RECT 4.1 1.455 4.33 3.315 ;
      RECT 2.305 1.455 4.1 1.685 ;
      RECT 3.4 3.085 4.1 3.315 ;
      RECT 3.17 3.085 3.4 3.685 ;
      RECT 3.06 3.345 3.17 3.685 ;
      RECT 2.075 1.075 2.305 1.685 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.23 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.39 2.185 3.82 2.72 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2626 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.58 2.265 3.085 2.785 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2914 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1554 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.66 0.76 2.13 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.3459 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2614 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.405 1.56 2.91 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2624 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.84 1.92 2.12 2.15 ;
      RECT 1.24 1.82 1.84 2.15 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.64 -0.4 4.62 0.4 ;
      RECT 3.3 -0.4 3.64 1.22 ;
      RECT 0.52 -0.4 3.3 0.4 ;
      RECT 0.18 -0.4 0.52 1.34 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.96 4.64 4.62 5.44 ;
      RECT 1.62 3.765 1.96 5.44 ;
      RECT 0.52 4.64 1.62 5.44 ;
      RECT 0.18 3.555 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.78 3.64 4.12 4.145 ;
      RECT 2.68 3.915 3.78 4.145 ;
      RECT 2.34 3.3 2.68 4.145 ;
      RECT 1.24 3.3 2.34 3.53 ;
      RECT 0.9 3.3 1.24 3.895 ;
  END
END AOI32XL

MACRO AOI32X4
  CLASS CORE ;
  FOREIGN AOI32X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI32XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.323 ;
  ANTENNAPARTIALMETALAREA 1.0174 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7312 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.31 1.82 6.46 3.22 ;
      RECT 6.08 1.5 6.31 3.22 ;
      RECT 5.775 1.5 6.08 1.73 ;
      RECT 5.415 2.74 6.08 3.08 ;
      RECT 5.435 1.39 5.775 1.73 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.3526 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4204 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.585 2.38 3.785 3.08 ;
      RECT 3.35 2.175 3.585 3.08 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.2932 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1501 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.12 2.38 2.63 2.955 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.3281 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.219 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.575 0.765 2.1 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.351 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.38 1.495 2.885 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2306 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.725 2.075 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.42 -0.4 6.6 0.4 ;
      RECT 6.08 -0.4 6.42 0.955 ;
      RECT 5.08 -0.4 6.08 0.4 ;
      RECT 4.85 -0.4 5.08 0.95 ;
      RECT 3.68 -0.4 4.85 0.4 ;
      RECT 3.34 -0.4 3.68 0.575 ;
      RECT 0.52 -0.4 3.34 0.4 ;
      RECT 0.18 -0.4 0.52 1.22 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.395 4.64 6.6 5.44 ;
      RECT 6.055 3.705 6.395 5.44 ;
      RECT 5.11 4.64 6.055 5.44 ;
      RECT 4.77 3.705 5.11 5.44 ;
      RECT 1.78 4.64 4.77 5.44 ;
      RECT 1.44 4.465 1.78 5.44 ;
      RECT 0.535 4.64 1.44 5.44 ;
      RECT 0.15 4.465 0.535 5.44 ;
      RECT 0 4.64 0.15 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.04 2.06 5.845 2.4 ;
      RECT 4.81 1.27 5.04 3.165 ;
      RECT 4.55 1.27 4.81 1.5 ;
      RECT 4.385 2.935 4.81 3.165 ;
      RECT 4.52 1.86 4.575 2.2 ;
      RECT 4.32 0.665 4.55 1.5 ;
      RECT 4.235 1.855 4.52 2.2 ;
      RECT 4.045 2.88 4.385 3.22 ;
      RECT 4.075 0.665 4.32 0.895 ;
      RECT 4.055 1.855 4.235 2.145 ;
      RECT 3.825 1.125 4.055 2.145 ;
      RECT 3.735 3.585 3.845 3.925 ;
      RECT 3.12 1.125 3.825 1.355 ;
      RECT 3.505 3.585 3.735 4.33 ;
      RECT 2.405 4.1 3.505 4.33 ;
      RECT 3.12 3.385 3.125 3.725 ;
      RECT 2.89 1.125 3.12 3.725 ;
      RECT 2.36 1.125 2.89 1.355 ;
      RECT 2.785 3.385 2.89 3.725 ;
      RECT 2.175 3.385 2.405 4.33 ;
      RECT 2.02 1.015 2.36 1.355 ;
      RECT 2.065 3.385 2.175 3.725 ;
      RECT 1.08 3.44 2.065 3.67 ;
      RECT 0.74 3.385 1.08 3.725 ;
  END
END AOI32X4

MACRO AOI32X2
  CLASS CORE ;
  FOREIGN AOI32X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI32XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.9958 ;
  ANTENNAPARTIALMETALAREA 2.2426 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.4145 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.815 1.46 7.045 3.315 ;
      RECT 6.74 1.46 6.815 1.845 ;
      RECT 6.375 3.085 6.815 3.315 ;
      RECT 6.27 1.46 6.74 1.69 ;
      RECT 6.035 3.03 6.375 3.37 ;
      RECT 6.04 1.18 6.27 1.69 ;
      RECT 3.245 1.18 6.04 1.41 ;
      RECT 5.095 3.075 6.035 3.305 ;
      RECT 4.755 3.02 5.095 3.36 ;
      RECT 3.015 0.795 3.245 1.41 ;
      RECT 2.02 0.795 3.015 1.025 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.6609 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2648 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.505 2.545 6.325 2.775 ;
      RECT 4.275 1.845 4.505 2.775 ;
      RECT 4.175 1.845 4.275 2.13 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.3169 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3939 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.32 1.82 5.8 2.13 ;
      RECT 4.98 1.82 5.32 2.31 ;
      RECT 4.975 1.82 4.98 2.13 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 0.9677 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.6693 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.605 2.39 3.835 2.905 ;
      RECT 3.44 2.63 3.605 2.905 ;
      RECT 0.645 2.675 3.44 2.905 ;
      RECT 0.415 2.405 0.645 2.905 ;
      RECT 0.215 2.405 0.415 2.635 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 0.6108 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.809 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.78 1.845 3.165 2.425 ;
      RECT 1.095 2.195 2.78 2.425 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 0.238 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3409 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.01 1.735 2.12 1.965 ;
      RECT 1.78 1.285 2.01 1.965 ;
      RECT 1.535 1.285 1.78 1.515 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.84 -0.4 7.26 0.4 ;
      RECT 6.5 -0.4 6.84 1.22 ;
      RECT 4.24 -0.4 6.5 0.4 ;
      RECT 3.9 -0.4 4.24 0.575 ;
      RECT 0.465 -0.4 3.9 0.4 ;
      RECT 0.235 -0.4 0.465 1.43 ;
      RECT 0 -0.4 0.235 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.725 4.64 7.26 5.44 ;
      RECT 3.385 4.09 3.725 5.44 ;
      RECT 2.445 4.64 3.385 5.44 ;
      RECT 2.105 4.09 2.445 5.44 ;
      RECT 1.16 4.64 2.105 5.44 ;
      RECT 0.82 4.09 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.675 3.765 7.015 4.105 ;
      RECT 5.735 3.82 6.675 4.05 ;
      RECT 5.395 3.765 5.735 4.105 ;
      RECT 4.455 3.82 5.395 4.05 ;
      RECT 4.345 3.765 4.455 4.105 ;
      RECT 4.115 3.41 4.345 4.105 ;
      RECT 3.085 3.41 4.115 3.64 ;
      RECT 2.745 3.355 3.085 3.695 ;
      RECT 1.805 3.4 2.745 3.63 ;
      RECT 1.465 3.345 1.805 3.685 ;
      RECT 0.52 3.4 1.465 3.63 ;
      RECT 0.18 3.345 0.52 3.685 ;
  END
END AOI32X2

MACRO AOI32X1
  CLASS CORE ;
  FOREIGN AOI32X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI32XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1584 ;
  ANTENNAPARTIALMETALAREA 1.3384 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.3706 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.175 0.935 4.405 3.445 ;
      RECT 4.1 0.935 4.175 1.285 ;
      RECT 3.06 3.215 4.175 3.445 ;
      RECT 2.02 0.935 4.1 1.165 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.2992 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.115 1.6 3.745 2.075 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.2142 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.53 2.35 3.16 2.69 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2772 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1448 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.68 0.8 2.1 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.2753 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1236 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.4 1.48 2.855 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3888 ;
  ANTENNAPARTIALMETALAREA 0.3234 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.219 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.61 2.12 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.71 -0.4 4.62 0.4 ;
      RECT 3.37 -0.4 3.71 0.575 ;
      RECT 0.465 -0.4 3.37 0.4 ;
      RECT 0.235 -0.4 0.465 1.43 ;
      RECT 0 -0.4 0.235 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.96 4.64 4.62 5.44 ;
      RECT 1.62 3.82 1.96 5.44 ;
      RECT 0.52 4.64 1.62 5.44 ;
      RECT 0.18 3.295 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.625 3.815 4.12 4.045 ;
      RECT 2.395 3.36 2.625 4.045 ;
      RECT 0.9 3.36 2.395 3.59 ;
  END
END AOI32X1

MACRO AOI31XL
  CLASS CORE ;
  FOREIGN AOI31XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.762 ;
  ANTENNAPARTIALMETALAREA 0.6876 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4026 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.065 1.175 3.085 1.515 ;
      RECT 2.835 1.175 3.065 3.32 ;
      RECT 2.02 1.175 2.835 1.405 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.2355 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0653 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.355 2.375 2.585 2.755 ;
      RECT 1.96 2.38 2.355 2.755 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2223 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.6 0.52 2.185 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.2397 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.38 1.485 2.73 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNAPARTIALMETALAREA 0.3415 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2773 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.54 1.64 2.28 2.1 ;
      RECT 1.535 1.845 1.54 2.075 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.065 -0.4 3.3 0.4 ;
      RECT 2.725 -0.4 3.065 0.575 ;
      RECT 0.52 -0.4 2.725 0.4 ;
      RECT 0.18 -0.4 0.52 1.22 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.84 4.64 3.3 5.44 ;
      RECT 1.5 4.465 1.84 5.44 ;
      RECT 0.545 4.64 1.5 5.44 ;
      RECT 0.175 4.465 0.545 5.44 ;
      RECT 0 4.64 0.175 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.74 3.19 2.4 3.53 ;
  END
END AOI31XL

MACRO AOI31X4
  CLASS CORE ;
  FOREIGN AOI31X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI31XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3334 ;
  ANTENNAPARTIALMETALAREA 0.9985 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.869 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.74 1.82 5.8 3.22 ;
      RECT 5.42 1.415 5.74 3.22 ;
      RECT 4.685 1.415 5.42 1.645 ;
      RECT 4.69 2.8 5.42 3.03 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2052 ;
  ANTENNAPARTIALMETALAREA 0.3049 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.625 1.8 3.16 2.37 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2185 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0123 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.525 0.52 2.1 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.3484 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2614 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.745 2.38 1.265 3.05 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2448 ;
  ANTENNAPARTIALMETALAREA 0.2132 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.415 1.72 1.935 2.13 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.67 -0.4 5.94 0.4 ;
      RECT 5.33 -0.4 5.67 0.96 ;
      RECT 4.385 -0.4 5.33 0.4 ;
      RECT 4.045 -0.4 4.385 0.96 ;
      RECT 2.96 -0.4 4.045 0.4 ;
      RECT 2.62 -0.4 2.96 0.575 ;
      RECT 0.52 -0.4 2.62 0.4 ;
      RECT 0.18 -0.4 0.52 1.29 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.615 4.64 5.94 5.44 ;
      RECT 5.385 3.735 5.615 5.44 ;
      RECT 4.385 4.64 5.385 5.44 ;
      RECT 4.045 3.76 4.385 5.44 ;
      RECT 1.64 4.64 4.045 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0.52 4.64 1.3 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.09 2.035 5.185 2.4 ;
      RECT 3.86 1.315 4.09 3.435 ;
      RECT 3.605 1.315 3.86 1.545 ;
      RECT 3.68 3.205 3.86 3.435 ;
      RECT 3.45 3.205 3.68 4.375 ;
      RECT 3.39 1.86 3.62 2.93 ;
      RECT 3.375 0.64 3.605 1.545 ;
      RECT 3.325 4.145 3.45 4.375 ;
      RECT 3.065 2.7 3.39 2.93 ;
      RECT 2.835 2.7 3.065 3.64 ;
      RECT 2.395 2.7 2.835 2.93 ;
      RECT 0.74 3.525 2.4 3.755 ;
      RECT 2.165 1.115 2.395 2.93 ;
      RECT 2.075 1.115 2.165 1.485 ;
  END
END AOI31X4

MACRO AOI31X2
  CLASS CORE ;
  FOREIGN AOI31X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI31XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5795 ;
  ANTENNAPARTIALMETALAREA 1.6848 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.9924 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.795 2.635 5.025 3.36 ;
      RECT 4.76 2.635 4.795 2.965 ;
      RECT 4.405 2.635 4.76 2.865 ;
      RECT 4.175 1.125 4.405 2.865 ;
      RECT 1.79 1.125 4.175 1.355 ;
      RECT 1.56 0.665 1.79 1.355 ;
      RECT 0.18 0.665 1.56 0.895 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6546 ;
  ANTENNAPARTIALMETALAREA 0.2833 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1289 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.635 1.82 5.18 2.34 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 0.4604 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2101 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.735 2.28 1.965 ;
      RECT 0.875 1.285 1.18 1.965 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 0.6132 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.16 2.215 3.275 2.445 ;
      RECT 2.78 1.845 3.16 2.445 ;
      RECT 1.22 2.215 2.78 2.445 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7842 ;
  ANTENNAPARTIALMETALAREA 1.1461 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.2735 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.675 2.06 3.905 2.905 ;
      RECT 0.52 2.675 3.675 2.905 ;
      RECT 0.14 2.31 0.52 2.905 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.96 -0.4 5.94 0.4 ;
      RECT 4.94 -0.4 4.96 0.575 ;
      RECT 4.71 -0.4 4.94 1.34 ;
      RECT 4.62 -0.4 4.71 0.575 ;
      RECT 2.36 -0.4 4.62 0.4 ;
      RECT 2.02 -0.4 2.36 0.895 ;
      RECT 0 -0.4 2.02 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.72 4.64 5.94 5.44 ;
      RECT 3.38 3.765 3.72 5.44 ;
      RECT 2.44 4.64 3.38 5.44 ;
      RECT 2.1 3.765 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 3.765 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.19 3.82 5.72 4.05 ;
      RECT 3.96 3.135 4.19 4.05 ;
      RECT 0.18 3.135 3.96 3.365 ;
  END
END AOI31X2

MACRO AOI31X1
  CLASS CORE ;
  FOREIGN AOI31X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI31XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.948 ;
  ANTENNAPARTIALMETALAREA 0.9721 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5633 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.025 0.845 3.085 3.175 ;
      RECT 2.855 0.845 3.025 4.025 ;
      RECT 2.78 0.845 2.855 1.54 ;
      RECT 2.795 2.945 2.855 4.025 ;
      RECT 2.02 0.845 2.78 1.075 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3273 ;
  ANTENNAPARTIALMETALAREA 0.249 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1236 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.62 2.105 2.625 2.45 ;
      RECT 2.23 2.105 2.62 2.66 ;
      RECT 2.12 2.38 2.23 2.66 ;
     END
  END B0

  PIN A2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3921 ;
  ANTENNAPARTIALMETALAREA 0.2413 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.765 0.52 2.4 ;
     END
  END A2

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3921 ;
  ANTENNAPARTIALMETALAREA 0.2277 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0123 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.345 1.295 2.805 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3921 ;
  ANTENNAPARTIALMETALAREA 0.2064 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 1.67 1.94 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.12 -0.4 3.3 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 0.52 -0.4 2.78 0.4 ;
      RECT 0.18 -0.4 0.52 0.895 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.8 4.64 3.3 5.44 ;
      RECT 1.46 3.78 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.785 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.82 3.04 2.44 3.27 ;
  END
END AOI31X1

MACRO AOI2BB2XL
  CLASS CORE ;
  FOREIGN AOI2BB2XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7588 ;
  ANTENNAPARTIALMETALAREA 0.7279 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5987 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.975 2.43 4.205 3.555 ;
      RECT 3.745 2.43 3.975 2.66 ;
      RECT 3.515 1.275 3.745 2.66 ;
      RECT 3.09 1.275 3.515 1.505 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2135 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.135 2.38 2.5 2.965 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2673 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1872 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.815 1.885 3.16 2.66 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.3136 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1925 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.59 0.755 2.1 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2755 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.495 1.18 3.22 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.1 -0.4 4.62 0.4 ;
      RECT 3.76 -0.4 4.1 0.575 ;
      RECT 2.12 -0.4 3.76 0.4 ;
      RECT 1.78 -0.4 2.12 0.575 ;
      RECT 0.52 -0.4 1.78 0.4 ;
      RECT 0.18 -0.4 0.52 1.22 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.78 4.64 4.62 5.44 ;
      RECT 2.44 4.465 2.78 5.44 ;
      RECT 0.52 4.64 2.44 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.975 0.81 4.205 2.095 ;
      RECT 1.64 0.81 3.975 1.04 ;
      RECT 3.2 3.635 3.54 3.975 ;
      RECT 2.165 3.69 3.2 3.92 ;
      RECT 1.935 3.215 2.165 3.92 ;
      RECT 1.41 0.81 1.64 4.28 ;
      RECT 0.98 0.99 1.41 1.22 ;
      RECT 1.395 3.92 1.41 4.28 ;
  END
END AOI2BB2XL

MACRO AOI2BB2X4
  CLASS CORE ;
  FOREIGN AOI2BB2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.9 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB2XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.3539 ;
  ANTENNAPARTIALMETALAREA 2.6832 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.7872 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.06 0.7 8.44 2.1 ;
      RECT 3.535 1.13 8.06 1.36 ;
      RECT 3.52 4.11 4.74 4.34 ;
      RECT 3.52 0.93 3.535 1.36 ;
      RECT 3.29 0.93 3.52 4.34 ;
      RECT 3.12 4.11 3.29 4.34 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 1.2344 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.9201 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.665 2.465 8.74 2.695 ;
      RECT 7.435 1.84 7.665 2.695 ;
      RECT 5.065 1.84 7.435 2.07 ;
      RECT 4.495 1.84 5.065 2.075 ;
      RECT 4.265 1.84 4.495 2.325 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.2146 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.955 2.38 6.46 2.805 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6048 ;
  ANTENNAPARTIALMETALAREA 1.3329 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.3494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.145 2.965 2.425 3.195 ;
      RECT 1.915 1.93 2.145 4.165 ;
      RECT 0.52 3.935 1.915 4.165 ;
      RECT 0.475 3.755 0.52 4.165 ;
      RECT 0.245 2.36 0.475 4.165 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6048 ;
  ANTENNAPARTIALMETALAREA 0.2326 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.75 1.715 1.22 2.21 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.095 -0.4 9.9 0.4 ;
      RECT 6.755 -0.4 7.095 0.895 ;
      RECT 4.31 -0.4 6.755 0.4 ;
      RECT 3.97 -0.4 4.31 0.895 ;
      RECT 2.485 -0.4 3.97 0.4 ;
      RECT 2.145 -0.4 2.485 0.575 ;
      RECT 0.915 -0.4 2.145 0.4 ;
      RECT 0.575 -0.4 0.915 0.895 ;
      RECT 0 -0.4 0.575 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.58 4.64 9.9 5.44 ;
      RECT 8.24 4.055 8.58 5.44 ;
      RECT 7.3 4.64 8.24 5.44 ;
      RECT 6.96 4.055 7.3 5.44 ;
      RECT 6.02 4.64 6.96 5.44 ;
      RECT 5.68 4.055 6.02 5.44 ;
      RECT 2.76 4.64 5.68 5.44 ;
      RECT 2.42 4.465 2.76 5.44 ;
      RECT 0.52 4.64 2.42 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.76 3.095 9.22 3.325 ;
      RECT 2.825 1.135 3.055 2.26 ;
      RECT 1.68 1.135 2.825 1.365 ;
      RECT 1.45 1.135 1.68 3.295 ;
      RECT 1.365 1.135 1.45 1.365 ;
      RECT 1.355 2.93 1.45 3.295 ;
  END
END AOI2BB2X4

MACRO AOI2BB2X2
  CLASS CORE ;
  FOREIGN AOI2BB2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB2XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4691 ;
  ANTENNAPARTIALMETALAREA 1.7682 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.1938 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.6 1.285 5.725 1.515 ;
      RECT 5.37 0.805 5.6 4.105 ;
      RECT 2.87 0.805 5.37 1.035 ;
      RECT 4.84 3.875 5.37 4.105 ;
      RECT 4.465 3.875 4.84 4.37 ;
      RECT 4.405 4.06 4.465 4.37 ;
      RECT 4.06 4.14 4.405 4.37 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.7994 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5775 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.1 2.28 4.46 3.095 ;
      RECT 1.9 2.865 4.1 3.095 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.6738 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2807 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.805 1.59 5.09 2.09 ;
      RECT 2.495 1.59 4.805 1.82 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3132 ;
  ANTENNAPARTIALMETALAREA 0.2655 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.275 1.63 1.84 2.1 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3132 ;
  ANTENNAPARTIALMETALAREA 0.3002 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.87 0.52 2.66 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.98 -0.4 5.94 0.4 ;
      RECT 3.64 -0.4 3.98 0.575 ;
      RECT 1.915 -0.4 3.64 0.4 ;
      RECT 1.575 -0.4 1.915 1.275 ;
      RECT 0.52 -0.4 1.575 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.72 4.64 5.94 5.44 ;
      RECT 5.38 4.465 5.72 5.44 ;
      RECT 3.12 4.64 5.38 5.44 ;
      RECT 2.78 4.085 3.12 5.44 ;
      RECT 1.84 4.64 2.78 5.44 ;
      RECT 1.5 4.085 1.84 5.44 ;
      RECT 0 4.64 1.5 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.14 3.395 5.04 3.625 ;
      RECT 1.025 2.4 3.68 2.63 ;
      RECT 0.795 1.21 1.025 3.31 ;
      RECT 0.18 3.08 0.795 3.31 ;
  END
END AOI2BB2X2

MACRO AOI2BB2X1
  CLASS CORE ;
  FOREIGN AOI2BB2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB2XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.9092 ;
  ANTENNAPARTIALMETALAREA 1.1404 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.9 1.115 4.13 4.405 ;
      RECT 2.7 1.115 3.9 1.345 ;
      RECT 3.515 2.38 3.9 2.66 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3633 ;
  ANTENNAPARTIALMETALAREA 0.2425 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.955 2.775 2.5 3.22 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3633 ;
  ANTENNAPARTIALMETALAREA 0.2288 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2985 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.855 2.25 3.085 2.635 ;
      RECT 2.62 2.25 2.855 2.48 ;
      RECT 2.39 2.105 2.62 2.48 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2237 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.19 1.82 0.475 2.605 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2134 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9805 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.795 2.25 1.235 2.735 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.8 -0.4 4.62 0.4 ;
      RECT 3.46 -0.4 3.8 0.575 ;
      RECT 1.72 -0.4 3.46 0.4 ;
      RECT 1.38 -0.4 1.72 0.575 ;
      RECT 0.52 -0.4 1.38 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.9 4.64 4.62 5.44 ;
      RECT 2.56 4.09 2.9 5.44 ;
      RECT 0.52 4.64 2.56 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.29 3.45 3.54 3.68 ;
      RECT 3.235 1.575 3.465 1.99 ;
      RECT 1.7 1.575 3.235 1.805 ;
      RECT 2.06 3.45 2.29 4.375 ;
      RECT 1.84 4.145 2.06 4.375 ;
      RECT 1.47 1.575 1.7 3.42 ;
      RECT 1.065 1.575 1.47 1.805 ;
      RECT 1.355 3.05 1.47 3.42 ;
      RECT 0.835 1.315 1.065 1.805 ;
  END
END AOI2BB2X1

MACRO AOI2BB1XL
  CLASS CORE ;
  FOREIGN AOI2BB1XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6562 ;
  ANTENNAPARTIALMETALAREA 0.7659 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7736 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.905 3.525 3.085 3.755 ;
      RECT 2.675 1.62 2.905 3.81 ;
      RECT 2.105 1.62 2.675 1.85 ;
      RECT 1.875 1.46 2.105 1.85 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.234 ;
  ANTENNAPARTIALMETALAREA 0.2695 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.67 1.95 3.22 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2118 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9964 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.54 2.26 1.105 2.635 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2331 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0335 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.175 2.895 0.73 3.315 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.27 -0.4 3.3 0.4 ;
      RECT 0.93 -0.4 1.27 0.575 ;
      RECT 0 -0.4 0.93 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.64 4.64 3.3 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0 4.64 1.3 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.18 2.085 2.41 3.785 ;
      RECT 1.64 2.085 2.18 2.315 ;
      RECT 0.18 3.555 2.18 3.785 ;
      RECT 1.41 1.315 1.64 2.315 ;
      RECT 0.45 1.315 1.41 1.545 ;
  END
END AOI2BB1XL

MACRO AOI2BB1X4
  CLASS CORE ;
  FOREIGN AOI2BB1X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB1XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.685 ;
  ANTENNAPARTIALMETALAREA 1.9333 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.0772 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.16 2.965 6.44 3.195 ;
      RECT 5.875 2.94 6.16 3.22 ;
      RECT 5.8 1.335 5.875 3.755 ;
      RECT 5.645 1.335 5.8 4.34 ;
      RECT 4.165 1.335 5.645 1.565 ;
      RECT 5.42 2.94 5.645 4.34 ;
      RECT 3.7 2.965 5.42 3.195 ;
      RECT 3.935 1.335 4.165 1.73 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3086 ;
  ANTENNAPARTIALMETALAREA 0.2769 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.85 1.82 3.24 2.53 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6156 ;
  ANTENNAPARTIALMETALAREA 1.1419 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.5067 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.385 1.845 2.425 2.075 ;
      RECT 2.155 1.845 2.385 3.735 ;
      RECT 0.475 3.505 2.155 3.735 ;
      RECT 0.245 2.38 0.475 3.735 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6156 ;
  ANTENNAPARTIALMETALAREA 0.2265 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2879 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.985 1.845 1.215 2.72 ;
      RECT 0.875 1.845 0.985 2.075 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.52 -0.4 7.26 0.4 ;
      RECT 6.18 -0.4 6.52 0.575 ;
      RECT 4.94 -0.4 6.18 0.4 ;
      RECT 4.6 -0.4 4.94 0.895 ;
      RECT 3.465 -0.4 4.6 0.4 ;
      RECT 3.125 -0.4 3.465 0.895 ;
      RECT 2.04 -0.4 3.125 0.4 ;
      RECT 1.7 -0.4 2.04 0.895 ;
      RECT 0 -0.4 1.7 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.185 4.64 7.26 5.44 ;
      RECT 4.955 4.025 5.185 5.44 ;
      RECT 2.76 4.64 4.955 5.44 ;
      RECT 2.42 4.465 2.76 5.44 ;
      RECT 0.52 4.64 2.42 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.185 1.925 5.415 2.645 ;
      RECT 3.7 2.415 5.185 2.645 ;
      RECT 3.47 1.36 3.7 2.645 ;
      RECT 1.675 1.36 3.47 1.59 ;
      RECT 1.445 1.36 1.675 3.195 ;
      RECT 0.975 1.36 1.445 1.59 ;
      RECT 1.3 2.965 1.445 3.195 ;
  END
END AOI2BB1X4

MACRO AOI2BB1X2
  CLASS CORE ;
  FOREIGN AOI2BB1X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB1XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.296 ;
  ANTENNAPARTIALMETALAREA 1.5906 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.8688 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.075 1.355 4.305 3.215 ;
      RECT 2.855 1.355 4.075 1.585 ;
      RECT 3.085 2.985 4.075 3.215 ;
      RECT 2.96 2.985 3.085 3.755 ;
      RECT 2.62 2.985 2.96 3.795 ;
      RECT 2.625 1.26 2.855 1.585 ;
      RECT 2.395 0.68 2.625 1.585 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.648 ;
  ANTENNAPARTIALMETALAREA 0.5635 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8408 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.585 1.845 3.815 2.68 ;
      RECT 2.385 1.845 3.585 2.075 ;
      RECT 2.155 1.845 2.385 2.26 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3132 ;
  ANTENNAPARTIALMETALAREA 0.2808 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.69 2.33 1.375 2.74 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3132 ;
  ANTENNAPARTIALMETALAREA 0.2106 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.26 0.53 1.8 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.44 -0.4 4.62 0.4 ;
      RECT 3.1 -0.4 3.44 0.575 ;
      RECT 1.96 -0.4 3.1 0.4 ;
      RECT 1.62 -0.4 1.96 0.895 ;
      RECT 0.52 -0.4 1.62 0.4 ;
      RECT 0.18 -0.4 0.52 0.895 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.24 4.64 4.62 5.44 ;
      RECT 3.9 3.55 4.24 5.44 ;
      RECT 1.64 4.64 3.9 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0 4.64 1.3 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.84 2.505 3.2 2.735 ;
      RECT 1.61 1.795 1.84 3.2 ;
      RECT 1.185 1.795 1.61 2.025 ;
      RECT 0.52 2.97 1.61 3.2 ;
      RECT 0.955 0.77 1.185 2.025 ;
      RECT 0.18 2.97 0.52 3.78 ;
  END
END AOI2BB1X2

MACRO AOI2BB1X1
  CLASS CORE ;
  FOREIGN AOI2BB1X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI2BB1XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8825 ;
  ANTENNAPARTIALMETALAREA 0.8866 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.3301 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.91 1.225 3.085 3.195 ;
      RECT 2.855 1.225 2.91 4.14 ;
      RECT 2.09 1.225 2.855 1.455 ;
      RECT 2.68 2.965 2.855 4.14 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3168 ;
  ANTENNAPARTIALMETALAREA 0.2761 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1395 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.96 2.795 1.965 3.195 ;
      RECT 1.315 2.795 1.96 3.22 ;
     END
  END B0

  PIN A1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.2142 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.55 1.78 1.18 2.12 ;
     END
  END A1N

  PIN A0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1548 ;
  ANTENNAPARTIALMETALAREA 0.3102 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1978 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.38 0.8 2.85 ;
     END
  END A0N

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.27 -0.4 3.3 0.4 ;
      RECT 0.93 -0.4 1.27 0.575 ;
      RECT 0 -0.4 0.93 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.64 4.64 3.3 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0 4.64 1.3 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.43 2.105 2.62 2.465 ;
      RECT 2.2 1.875 2.43 3.755 ;
      RECT 1.695 1.875 2.2 2.105 ;
      RECT 0.18 3.525 2.2 3.755 ;
      RECT 1.465 1.305 1.695 2.105 ;
      RECT 0.45 1.305 1.465 1.535 ;
  END
END AOI2BB1X1

MACRO AOI22XL
  CLASS CORE ;
  FOREIGN AOI22XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.756 ;
  ANTENNAPARTIALMETALAREA 1.1172 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.247 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.93 1.185 3.16 3.425 ;
      RECT 2.855 1.185 2.93 1.515 ;
      RECT 2.44 3.195 2.93 3.425 ;
      RECT 1.84 1.185 2.855 1.415 ;
      RECT 2.1 3.14 2.44 3.48 ;
      RECT 1.5 1.13 1.84 1.47 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2304 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.665 0.62 2.145 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.262 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.19 2.35 1.53 2.725 ;
      RECT 0.8 2.38 1.19 2.725 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2258 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.625 2.4 2.68 2.74 ;
      RECT 2.08 2.36 2.625 2.74 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2384 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.205 1.785 2.21 2.1 ;
      RECT 1.765 1.73 2.205 2.1 ;
      RECT 1.53 1.785 1.765 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.08 -0.4 3.3 0.4 ;
      RECT 2.74 -0.4 3.08 0.575 ;
      RECT 0.52 -0.4 2.74 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.645 4.64 3.3 5.44 ;
      RECT 0.23 4.465 0.645 5.44 ;
      RECT 0 4.64 0.23 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.66 4.175 3.01 4.405 ;
      RECT 1.43 3.2 1.66 4.405 ;
      RECT 0.52 3.2 1.43 3.43 ;
      RECT 0.18 3.145 0.52 3.485 ;
  END
END AOI22XL

MACRO AOI22X4
  CLASS CORE ;
  FOREIGN AOI22X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.24 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI22XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 4.1709 ;
  ANTENNAPARTIALMETALAREA 3.8281 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 16.3293 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.44 1.845 8.67 4.135 ;
      RECT 8.365 1.26 8.44 2.66 ;
      RECT 7.48 3.905 8.44 4.135 ;
      RECT 8.06 1.205 8.365 2.66 ;
      RECT 0.18 1.205 8.06 1.435 ;
      RECT 7.165 3.905 7.48 4.34 ;
      RECT 7.04 4.06 7.165 4.34 ;
      RECT 4.66 4.11 7.04 4.34 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.7187 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5563 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.94 1.84 3.995 2.07 ;
      RECT 3.71 1.84 3.94 2.075 ;
      RECT 0.875 1.845 3.71 2.075 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.5715 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8779 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.425 2.465 2.845 2.695 ;
      RECT 2.195 2.405 2.425 2.695 ;
      RECT 0.42 2.465 2.195 2.695 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.742 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6464 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.76 1.845 6.92 2.075 ;
      RECT 4.61 1.845 4.76 2.1 ;
      RECT 4.38 1.845 4.61 2.745 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.4058 ;
  ANTENNAPARTIALMETALAREA 0.6911 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4291 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.55 2.115 7.78 2.635 ;
      RECT 5.065 2.405 7.55 2.635 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.92 -0.4 9.24 0.4 ;
      RECT 6.58 -0.4 6.92 0.915 ;
      RECT 4.36 -0.4 6.58 0.4 ;
      RECT 4.02 -0.4 4.36 0.915 ;
      RECT 1.8 -0.4 4.02 0.4 ;
      RECT 1.46 -0.4 1.8 0.915 ;
      RECT 0 -0.4 1.46 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.72 4.64 9.24 5.44 ;
      RECT 3.38 4.055 3.72 5.44 ;
      RECT 2.44 4.64 3.38 5.44 ;
      RECT 2.1 4.055 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 4.055 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.18 3.095 8.2 3.325 ;
  END
END AOI22X4

MACRO AOI22X2
  CLASS CORE ;
  FOREIGN AOI22X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI22XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.0062 ;
  ANTENNAPARTIALMETALAREA 1.8498 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.7609 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.495 1.35 5.725 3.195 ;
      RECT 1.46 1.35 5.495 1.58 ;
      RECT 5.08 2.965 5.495 3.195 ;
      RECT 4.835 2.965 5.08 3.315 ;
      RECT 3.46 3.085 4.835 3.315 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.6708 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2012 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.425 1.915 2.655 2.415 ;
      RECT 1.105 1.915 2.425 2.145 ;
      RECT 0.915 1.845 1.105 2.145 ;
      RECT 0.685 1.845 0.915 2.36 ;
      RECT 0.42 2.07 0.685 2.36 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.2071 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9805 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.22 2.405 1.765 2.785 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.6808 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3761 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.035 1.84 5.265 2.315 ;
      RECT 3.745 1.84 5.035 2.07 ;
      RECT 3.505 1.84 3.745 2.075 ;
      RECT 3.275 1.84 3.505 2.79 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.2133 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9911 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.94 2.38 4.48 2.775 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.36 -0.4 5.94 0.4 ;
      RECT 5.02 -0.4 5.36 0.575 ;
      RECT 2.92 -0.4 5.02 0.4 ;
      RECT 2.58 -0.4 2.92 0.575 ;
      RECT 0.52 -0.4 2.58 0.4 ;
      RECT 0.18 -0.4 0.52 1.345 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.44 4.64 5.94 5.44 ;
      RECT 2.1 3.665 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 3.665 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.025 3.72 5.72 3.95 ;
      RECT 3.025 3.075 3.08 3.305 ;
      RECT 2.795 3.075 3.025 3.95 ;
      RECT 0.18 3.075 2.795 3.305 ;
  END
END AOI22X2

MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI22XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.9772 ;
  ANTENNAPARTIALMETALAREA 1.0788 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.0456 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.93 1.115 3.16 3.165 ;
      RECT 2.855 1.115 2.93 1.515 ;
      RECT 2.48 2.935 2.93 3.165 ;
      RECT 1.8 1.115 2.855 1.345 ;
      RECT 2.14 2.935 2.48 3.275 ;
      RECT 1.46 1.06 1.8 1.4 ;
     END
  END Y

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.2397 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.19 1.77 0.53 2.475 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.2612 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.38 1.52 2.785 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3642 ;
  ANTENNAPARTIALMETALAREA 0.2259 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.115 2.26 2.68 2.66 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3642 ;
  ANTENNAPARTIALMETALAREA 0.2181 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1183 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.83 1.655 2.17 1.995 ;
      RECT 1.765 1.71 1.83 1.995 ;
      RECT 1.535 1.71 1.765 2.075 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.12 -0.4 3.3 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 0.52 -0.4 2.78 0.4 ;
      RECT 0.18 -0.4 0.52 1.45 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 3.3 5.44 ;
      RECT 0.84 4.465 1.18 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.78 3.585 3.12 3.925 ;
      RECT 1.84 3.695 2.78 3.925 ;
      RECT 1.5 3.635 1.84 3.975 ;
      RECT 0.52 3.69 1.5 3.92 ;
      RECT 0.18 3.05 0.52 3.92 ;
  END
END AOI22X1

MACRO AOI222XL
  CLASS CORE ;
  FOREIGN AOI222XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1848 ;
  ANTENNAPARTIALMETALAREA 1.7388 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.1779 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.835 1.135 5.065 3.095 ;
      RECT 0.18 1.135 4.835 1.365 ;
      RECT 4.76 2.635 4.835 3.095 ;
      RECT 3.965 2.865 4.76 3.095 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.235 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.385 1.27 2.885 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.52 2.37 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.2062 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9805 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.525 1.725 2.075 2.1 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.595 1.82 3.145 2.2 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.2432 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.17 1.845 4.52 2.54 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2736 ;
  ANTENNAPARTIALMETALAREA 0.209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.475 1.645 3.855 2.195 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.85 -0.4 5.28 0.4 ;
      RECT 4.51 -0.4 4.85 0.575 ;
      RECT 1.885 -0.4 4.51 0.4 ;
      RECT 1.545 -0.4 1.885 0.905 ;
      RECT 0 -0.4 1.545 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.16 4.64 5.28 5.44 ;
      RECT 0.82 4.41 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.08 4.145 4.865 4.375 ;
      RECT 0.74 3.365 2.98 3.595 ;
  END
END AOI222XL

MACRO AOI222X4
  CLASS CORE ;
  FOREIGN AOI222X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.92 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI222XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2895 ;
  ANTENNAPARTIALMETALAREA 0.9359 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5298 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.07 2.38 7.12 3.78 ;
      RECT 6.84 1.41 7.07 3.78 ;
      RECT 6.74 1.41 6.84 1.85 ;
      RECT 6.74 2.38 6.84 3.78 ;
      RECT 6.5 1.41 6.74 1.64 ;
      RECT 6.5 2.775 6.74 3.115 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.304 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.52 2.62 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.3243 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.87 1.605 1.56 2.075 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2035 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1819 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.535 2.405 2.42 2.635 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2755 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.78 2.12 3.16 2.845 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2413 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.125 2.2 4.48 2.88 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2527 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.44 1.67 3.82 2.335 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.48 -0.4 7.92 0.4 ;
      RECT 7.14 -0.4 7.48 0.955 ;
      RECT 6.16 -0.4 7.14 0.4 ;
      RECT 5.82 -0.4 6.16 0.955 ;
      RECT 4.74 -0.4 5.82 0.4 ;
      RECT 4.4 -0.4 4.74 0.575 ;
      RECT 2.5 -0.4 4.4 0.4 ;
      RECT 2.16 -0.4 2.5 0.575 ;
      RECT 0.68 -0.4 2.16 0.4 ;
      RECT 0.52 -0.4 0.68 0.41 ;
      RECT 0.18 -0.4 0.52 1.22 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.48 4.64 7.92 5.44 ;
      RECT 7.14 4.06 7.48 5.44 ;
      RECT 6.2 4.64 7.14 5.44 ;
      RECT 5.86 3.75 6.2 5.44 ;
      RECT 1.64 4.64 5.86 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0.52 4.64 1.3 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.015 2.225 6.505 2.455 ;
      RECT 5.785 1.205 6.015 2.96 ;
      RECT 5.1 1.205 5.785 1.435 ;
      RECT 5.425 2.73 5.785 2.96 ;
      RECT 4.94 2.185 5.47 2.415 ;
      RECT 5.195 2.73 5.425 3.11 ;
      RECT 4.71 1.695 4.94 3.5 ;
      RECT 2 4.18 4.78 4.41 ;
      RECT 4.295 1.695 4.71 1.925 ;
      RECT 3.88 3.27 4.71 3.5 ;
      RECT 4.065 1.115 4.295 1.925 ;
      RECT 3.63 1.115 4.065 1.345 ;
      RECT 3.28 0.99 3.63 1.345 ;
      RECT 1.46 0.99 3.28 1.22 ;
      RECT 0.74 3.41 2.9 3.64 ;
  END
END AOI222X4

MACRO AOI222X2
  CLASS CORE ;
  FOREIGN AOI222X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.24 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI222XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.4934 ;
  ANTENNAPARTIALMETALAREA 2.7079 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 12.3278 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.635 1.125 8.865 3.12 ;
      RECT 8.365 1.125 8.635 1.54 ;
      RECT 8.365 2.89 8.635 3.12 ;
      RECT 7.48 1.125 8.365 1.355 ;
      RECT 8.135 2.89 8.365 3.195 ;
      RECT 6.64 2.89 8.135 3.12 ;
      RECT 7.04 1.045 7.48 1.355 ;
      RECT 4.87 1.125 7.04 1.355 ;
      RECT 4.4 1.045 4.87 1.355 ;
      RECT 1.46 1.125 4.4 1.355 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.6168 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9892 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.32 2.335 2.68 2.605 ;
      RECT 1.105 2.375 2.32 2.605 ;
      RECT 0.575 2.375 1.105 2.635 ;
      RECT 0.345 2.19 0.575 2.635 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.3358 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2614 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.67 1.91 2.13 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.5163 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6235 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.515 1.845 5.76 2.075 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.216 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.175 2.345 4.92 2.635 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.5658 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8514 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.17 1.845 8.4 2.29 ;
      RECT 6.155 1.845 8.17 2.075 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.2235 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.705 2.335 7.45 2.635 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.695 -0.4 9.24 0.4 ;
      RECT 8.355 -0.4 8.695 0.895 ;
      RECT 6.13 -0.4 8.355 0.4 ;
      RECT 5.79 -0.4 6.13 0.895 ;
      RECT 3.23 -0.4 5.79 0.4 ;
      RECT 2.89 -0.4 3.23 0.895 ;
      RECT 0.52 -0.4 2.89 0.4 ;
      RECT 0.18 -0.4 0.52 1.22 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.08 4.64 9.24 5.44 ;
      RECT 2.74 3.765 3.08 5.44 ;
      RECT 1.8 4.64 2.74 5.44 ;
      RECT 1.46 3.765 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.765 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.44 3.82 8.9 4.05 ;
      RECT 0.82 2.89 5.7 3.12 ;
  END
END AOI222X2

MACRO AOI222X1
  CLASS CORE ;
  FOREIGN AOI222X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.28 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI222XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4547 ;
  ANTENNAPARTIALMETALAREA 1.6893 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.0295 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.835 1.18 5.065 3.12 ;
      RECT 0.18 1.18 4.835 1.41 ;
      RECT 4.085 2.89 4.835 3.12 ;
     END
  END Y

  PIN C1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2408 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 1.7 1.435 2.13 ;
     END
  END C1

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2608 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2031 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.845 0.46 2.66 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2588 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2561 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.84 2.125 2.21 2.635 ;
      RECT 1.535 2.405 1.84 2.635 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2189 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9964 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.645 1.82 3.16 2.245 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2451 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.1 1.82 4.48 2.465 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3993 ;
  ANTENNAPARTIALMETALAREA 0.2926 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.219 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.44 1.865 3.82 2.635 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.785 -0.4 5.28 0.4 ;
      RECT 4.445 -0.4 4.785 0.575 ;
      RECT 1.915 -0.4 4.445 0.4 ;
      RECT 1.575 -0.4 1.915 0.575 ;
      RECT 0 -0.4 1.575 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.8 4.64 5.28 5.44 ;
      RECT 1.46 3.79 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.89 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.165 3.82 5.065 4.05 ;
      RECT 2.665 2.875 3.145 3.105 ;
      RECT 2.435 2.875 2.665 3.43 ;
      RECT 0.82 3.2 2.435 3.43 ;
  END
END AOI222X1

MACRO AOI221XL
  CLASS CORE ;
  FOREIGN AOI221XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.9861 ;
  ANTENNAPARTIALMETALAREA 1.273 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.0261 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.175 0.99 4.405 3.12 ;
      RECT 4.1 0.99 4.175 1.285 ;
      RECT 3.88 2.89 4.175 3.12 ;
      RECT 2.175 0.99 4.1 1.22 ;
      RECT 1.945 0.675 2.175 1.22 ;
      RECT 1.765 0.675 1.945 0.98 ;
      RECT 1.46 0.675 1.765 0.905 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2556 ;
  ANTENNAPARTIALMETALAREA 0.2162 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.62 2.405 3.745 2.635 ;
      RECT 3.39 1.82 3.62 2.635 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.2983 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.315 0.52 2.1 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.2484 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.36 1.34 2.82 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.2626 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.565 1.57 3.085 2.075 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2808 ;
  ANTENNAPARTIALMETALAREA 0.2138 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2296 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.735 1.845 1.965 2.575 ;
      RECT 1.535 1.845 1.735 2.075 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.12 -0.4 4.62 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 0.52 -0.4 2.78 0.4 ;
      RECT 0.18 -0.4 0.52 0.895 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.64 4.64 4.62 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0.52 4.64 1.3 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2 4.18 3.46 4.41 ;
      RECT 2.56 2.82 2.9 3.64 ;
      RECT 1.08 3.41 2.56 3.64 ;
      RECT 0.74 3.11 1.08 3.93 ;
  END
END AOI221XL

MACRO AOI221X4
  CLASS CORE ;
  FOREIGN AOI221X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI221XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5876 ;
  ANTENNAPARTIALMETALAREA 1.0467 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6782 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.31 1.26 6.46 2.66 ;
      RECT 6.08 1.26 6.31 4.05 ;
      RECT 5.9 1.26 6.08 1.49 ;
      RECT 5.96 2.77 6.08 4.05 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.3136 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1925 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.13 1.565 3.745 2.075 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2717 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.94 0.52 2.655 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2363 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0918 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.51 1.22 3.195 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2304 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2561 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.655 2.38 3.085 2.635 ;
      RECT 2.425 2.11 2.655 2.635 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2571 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.535 1.82 1.94 2.455 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.92 -0.4 7.26 0.4 ;
      RECT 6.69 -0.4 6.92 1.58 ;
      RECT 5.52 -0.4 6.69 0.4 ;
      RECT 5.18 -0.4 5.52 0.895 ;
      RECT 3.12 -0.4 5.18 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 0.52 -0.4 2.78 0.4 ;
      RECT 0.18 -0.4 0.52 1.285 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.02 4.64 7.26 5.44 ;
      RECT 6.68 3.15 7.02 5.44 ;
      RECT 5.58 4.64 6.68 5.44 ;
      RECT 5.24 3.15 5.58 5.44 ;
      RECT 1.64 4.64 5.24 5.44 ;
      RECT 1.3 4.465 1.64 5.44 ;
      RECT 0.52 4.64 1.3 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.07 2.135 5.71 2.365 ;
      RECT 4.86 1.45 5.07 2.705 ;
      RECT 4.84 1.45 4.86 4.1 ;
      RECT 4.74 1.45 4.84 1.68 ;
      RECT 4.63 2.475 4.84 4.1 ;
      RECT 4.51 1.15 4.74 1.68 ;
      RECT 4.52 3.76 4.63 4.1 ;
      RECT 4.28 1.965 4.61 2.195 ;
      RECT 4.05 0.99 4.28 3.4 ;
      RECT 2.415 0.99 4.05 1.22 ;
      RECT 3.935 3.035 4.05 3.4 ;
      RECT 0.74 3.495 2.9 3.725 ;
      RECT 2.185 0.99 2.415 1.285 ;
      RECT 1.46 1.055 2.185 1.285 ;
  END
END AOI221X4

MACRO AOI221X2
  CLASS CORE ;
  FOREIGN AOI221X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.92 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI221XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.9726 ;
  ANTENNAPARTIALMETALAREA 1.8936 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.8245 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.815 1.31 7.045 3.51 ;
      RECT 5.495 1.31 6.815 1.54 ;
      RECT 6.64 3.17 6.815 3.51 ;
      RECT 5.245 1.26 5.495 1.54 ;
      RECT 5.015 0.945 5.245 1.54 ;
      RECT 1.46 0.945 5.015 1.175 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7284 ;
  ANTENNAPARTIALMETALAREA 0.2921 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.59 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.33 1.845 6.56 2.28 ;
      RECT 5.495 1.845 6.33 2.075 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8004 ;
  ANTENNAPARTIALMETALAREA 0.6698 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0899 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.5 2.07 2.68 2.345 ;
      RECT 2.12 1.82 2.5 2.345 ;
      RECT 0.29 2.115 2.12 2.345 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8004 ;
  ANTENNAPARTIALMETALAREA 0.285 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.575 1.56 1.805 ;
      RECT 0.8 1.285 1.18 1.805 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8004 ;
  ANTENNAPARTIALMETALAREA 0.5899 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9627 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.745 2.5 5.93 2.73 ;
      RECT 3.515 2.405 3.745 2.73 ;
      RECT 3.46 2.5 3.515 2.73 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.8004 ;
  ANTENNAPARTIALMETALAREA 0.2392 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0441 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.1 1.665 4.65 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.17 -0.4 7.92 0.4 ;
      RECT 5.83 -0.4 6.17 0.895 ;
      RECT 3.28 -0.4 5.83 0.4 ;
      RECT 2.94 -0.4 3.28 0.575 ;
      RECT 0.52 -0.4 2.94 0.4 ;
      RECT 0.18 -0.4 0.52 0.895 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.08 4.64 7.92 5.44 ;
      RECT 2.74 3.73 3.08 5.44 ;
      RECT 1.8 4.64 2.74 5.44 ;
      RECT 1.46 3.73 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.73 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.44 4.04 7.62 4.27 ;
      RECT 3.56 3.225 5.7 3.455 ;
      RECT 3.33 2.97 3.56 3.455 ;
      RECT 0.82 2.97 3.33 3.2 ;
  END
END AOI221X2

MACRO AOI221X1
  CLASS CORE ;
  FOREIGN AOI221X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI221XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3164 ;
  ANTENNAPARTIALMETALAREA 1.1981 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.7028 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.175 1.08 4.405 3.195 ;
      RECT 2.5 1.08 4.175 1.31 ;
      RECT 4.14 2.635 4.175 3.165 ;
      RECT 2.475 0.955 2.5 1.31 ;
      RECT 2.245 0.795 2.475 1.31 ;
      RECT 1.46 0.795 2.245 1.025 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3646 ;
  ANTENNAPARTIALMETALAREA 0.2346 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.325 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.71 2.405 3.745 2.635 ;
      RECT 3.48 1.65 3.71 2.635 ;
     END
  END C0

  PIN B1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4006 ;
  ANTENNAPARTIALMETALAREA 0.2242 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.175 1.285 0.52 1.935 ;
     END
  END B1

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4006 ;
  ANTENNAPARTIALMETALAREA 0.2612 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.185 1.35 2.66 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4006 ;
  ANTENNAPARTIALMETALAREA 0.2231 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.272 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.855 1.59 3.085 2.075 ;
      RECT 2.37 1.59 2.855 1.82 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4006 ;
  ANTENNAPARTIALMETALAREA 0.2389 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.535 1.285 1.99 1.81 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.12 -0.4 4.62 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 0.52 -0.4 2.78 0.4 ;
      RECT 0.18 -0.4 0.52 1.025 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.8 4.64 4.62 5.44 ;
      RECT 1.46 3.785 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 3.785 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.165 3.62 3.785 3.85 ;
      RECT 0.82 2.895 3.145 3.125 ;
  END
END AOI221X1

MACRO AOI21XL
  CLASS CORE ;
  FOREIGN AOI21XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.679 ;
  ANTENNAPARTIALMETALAREA 0.6934 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4397 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.39 1.24 2.425 2.635 ;
      RECT 2.195 1.24 2.39 3.485 ;
      RECT 1.46 1.24 2.195 1.47 ;
      RECT 2.16 2.405 2.195 3.485 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.2137 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0017 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.365 1.725 1.935 2.1 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2135 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.17 1.75 0.52 2.36 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.252 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0918 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.38 1.43 2.78 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.36 -0.4 2.64 0.4 ;
      RECT 2.02 -0.4 2.36 0.575 ;
      RECT 0.52 -0.4 2.02 0.4 ;
      RECT 0.18 -0.4 0.52 1.455 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 4.64 2.64 5.44 ;
      RECT 0.84 4.465 1.18 5.44 ;
      RECT 0 4.64 0.84 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.64 4.18 1.88 4.41 ;
      RECT 1.41 4 1.64 4.41 ;
      RECT 0.465 4 1.41 4.23 ;
      RECT 0.235 3.145 0.465 4.23 ;
  END
END AOI21XL

MACRO AOI21X4
  CLASS CORE ;
  FOREIGN AOI21X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI21XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.904 ;
  ANTENNAPARTIALMETALAREA 2.6215 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.1777 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.115 3.765 6.28 4.105 ;
      RECT 5.94 2.43 6.115 4.105 ;
      RECT 5.885 2.43 5.94 4.05 ;
      RECT 5.8 2.43 5.885 2.66 ;
      RECT 5 3.82 5.885 4.05 ;
      RECT 5.42 1.26 5.8 2.66 ;
      RECT 4.835 1.415 5.42 1.645 ;
      RECT 4.66 3.765 5 4.105 ;
      RECT 4.43 1.15 4.835 1.645 ;
      RECT 0.18 1.15 4.43 1.38 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.2594 ;
  ANTENNAPARTIALMETALAREA 0.348 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.54 2.085 5.14 2.665 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.8876 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6146 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.915 1.9 4.025 2.24 ;
      RECT 3.685 1.645 3.915 2.24 ;
      RECT 2.425 1.645 3.685 1.875 ;
      RECT 1.805 1.645 2.425 2.075 ;
      RECT 1.52 1.645 1.805 2.13 ;
      RECT 1.465 1.79 1.52 2.13 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.449 ;
  ANTENNAPARTIALMETALAREA 0.7757 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.71 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.96 2.405 3.085 2.635 ;
      RECT 2.73 2.225 2.96 2.635 ;
      RECT 0.8 2.395 2.73 2.625 ;
      RECT 0.76 2.38 0.8 2.625 ;
      RECT 0.53 1.97 0.76 2.625 ;
      RECT 0.42 1.97 0.53 2.41 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.685 -0.4 6.6 0.4 ;
      RECT 5.345 -0.4 5.685 0.575 ;
      RECT 4.365 -0.4 5.345 0.4 ;
      RECT 4.025 -0.4 4.365 0.895 ;
      RECT 1.805 -0.4 4.025 0.4 ;
      RECT 1.465 -0.4 1.805 0.895 ;
      RECT 0 -0.4 1.465 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.72 4.64 6.6 5.44 ;
      RECT 3.38 3.89 3.72 5.44 ;
      RECT 2.44 4.64 3.38 5.44 ;
      RECT 2.1 3.89 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 3.89 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.18 2.93 5.64 3.16 ;
  END
END AOI21X4

MACRO AOI21X2
  CLASS CORE ;
  FOREIGN AOI21X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.62 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI21XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5635 ;
  ANTENNAPARTIALMETALAREA 1.49 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.8105 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.66 1.45 3.89 3.315 ;
      RECT 3.08 1.45 3.66 1.68 ;
      RECT 3.515 2.965 3.66 3.315 ;
      RECT 3.46 3.085 3.515 3.315 ;
      RECT 2.74 1.125 3.08 1.68 ;
      RECT 1.065 1.45 2.74 1.68 ;
      RECT 0.835 1.235 1.065 1.68 ;
      RECT 0.52 1.235 0.835 1.465 ;
      RECT 0.18 1.125 0.52 1.465 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6546 ;
  ANTENNAPARTIALMETALAREA 0.2468 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1342 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.95 2.035 3.325 2.635 ;
      RECT 2.855 2.405 2.95 2.635 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.321 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4522 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.5 1.84 2.81 ;
      RECT 0.875 2.405 1.105 2.81 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7266 ;
  ANTENNAPARTIALMETALAREA 0.6576 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1535 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 1.92 2.71 2.15 ;
      RECT 0.14 1.82 0.52 2.225 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.845 -0.4 4.62 0.4 ;
      RECT 3.505 -0.4 3.845 0.575 ;
      RECT 1.8 -0.4 3.505 0.4 ;
      RECT 1.46 -0.4 1.8 1.22 ;
      RECT 0 -0.4 1.46 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.44 4.64 4.62 5.44 ;
      RECT 2.1 3.665 2.44 5.44 ;
      RECT 1.16 4.64 2.1 5.44 ;
      RECT 0.82 3.665 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.1 3.665 4.44 4.005 ;
      RECT 3.095 3.665 4.1 3.895 ;
      RECT 2.865 3.075 3.095 3.895 ;
      RECT 0.18 3.075 2.865 3.305 ;
  END
END AOI21X2

MACRO AOI21X1
  CLASS CORE ;
  FOREIGN AOI21X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI21XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8992 ;
  ANTENNAPARTIALMETALAREA 0.9339 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1658 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.275 1.35 2.505 3.95 ;
      RECT 1.8 1.35 2.275 1.58 ;
      RECT 2.195 2.965 2.275 3.95 ;
      RECT 2.1 3.61 2.195 3.95 ;
      RECT 1.46 1.24 1.8 1.58 ;
     END
  END Y

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3282 ;
  ANTENNAPARTIALMETALAREA 0.2545 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.378 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.8 1.845 2.045 2.635 ;
      RECT 1.535 1.845 1.8 2.075 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3642 ;
  ANTENNAPARTIALMETALAREA 0.2576 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 2.065 0.53 2.585 ;
      RECT 0.19 1.82 0.52 2.585 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3642 ;
  ANTENNAPARTIALMETALAREA 0.3806 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.9981 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.385 1.43 2.615 ;
      RECT 0.875 1.285 1.105 2.615 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.36 -0.4 2.64 0.4 ;
      RECT 2.02 -0.4 2.36 0.575 ;
      RECT 0.52 -0.4 2.02 0.4 ;
      RECT 0.18 -0.4 0.52 1.465 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.16 4.64 2.64 5.44 ;
      RECT 0.82 3.515 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.18 2.925 1.8 3.155 ;
  END
END AOI21X1

MACRO NAND2X0_LVT
  CLASS CORE ;
  FOREIGN NAND2X0_LVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5216 ;
  ANTENNAPARTIALMETALAREA 0.7362 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3549 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.705 3.19 3.82 3.78 ;
      RECT 3.475 1.015 3.705 3.78 ;
      RECT 3.42 3.19 3.475 3.78 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1584 ;
  ANTENNAPARTIALMETALAREA 0.274 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.54 2.405 3.105 2.89 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1584 ;
  ANTENNAPARTIALMETALAREA 0.2869 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2031 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.135 1.84 2.89 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1584 ;
  ANTENNAPARTIALMETALAREA 0.2869 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2031 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.135 1.18 2.89 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1584 ;
  ANTENNAPARTIALMETALAREA 0.2565 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1183 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.545 0.52 3.22 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3 -0.4 3.96 0.4 ;
      RECT 2.66 -0.4 3 0.575 ;
      RECT 0 -0.4 2.66 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.1 4.64 3.96 5.44 ;
      RECT 0.93 4.465 3.1 5.44 ;
      RECT 0 4.64 0.93 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.3 1.54 3.225 1.91 ;
      RECT 2.26 0.975 2.3 3.46 ;
      RECT 2.07 0.975 2.26 3.725 ;
      RECT 0.52 0.975 2.07 1.205 ;
      RECT 1.92 3.155 2.07 3.725 ;
      RECT 0.52 3.495 1.92 3.725 ;
      RECT 0.18 0.975 0.52 1.315 ;
  END
END NAND2X0_LVT

MACRO AND4X4
  CLASS CORE ;
  FOREIGN AND4X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ NAND2X0_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.6126 ;
  ANTENNAPARTIALMETALAREA 1.4405 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.876 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.385 2.38 6.46 3.78 ;
      RECT 6.155 1.495 6.385 3.78 ;
      RECT 6.085 1.39 6.155 3.78 ;
      RECT 6.08 1.39 6.085 1.845 ;
      RECT 6.08 2.38 6.085 3.78 ;
      RECT 5.7 1.39 6.08 1.73 ;
      RECT 5.56 3.425 6.08 3.78 ;
      RECT 5.22 3.425 5.56 4.365 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5202 ;
  ANTENNAPARTIALMETALAREA 1.7445 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.9606 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.82 1.845 4.95 2.075 ;
      RECT 4.59 1.845 4.82 2.73 ;
      RECT 4.405 2.38 4.59 2.73 ;
      RECT 4.275 2.5 4.405 2.73 ;
      RECT 4.045 2.5 4.275 3.73 ;
      RECT 0.525 3.5 4.045 3.73 ;
      RECT 0.525 2.69 0.53 3.22 ;
      RECT 0.295 2.69 0.525 3.73 ;
      RECT 0.14 2.69 0.295 3.22 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5202 ;
  ANTENNAPARTIALMETALAREA 1.2806 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.6975 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.585 1.59 3.815 3.03 ;
      RECT 3.44 1.59 3.585 1.845 ;
      RECT 1.25 1.59 3.44 1.82 ;
      RECT 1.25 2.265 1.32 2.67 ;
      RECT 1.02 1.59 1.25 2.67 ;
      RECT 0.8 2.07 1.02 2.67 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5202 ;
  ANTENNAPARTIALMETALAREA 0.4775 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.1995 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.78 2.055 3.16 2.64 ;
      RECT 1.67 2.055 2.78 2.285 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5202 ;
  ANTENNAPARTIALMETALAREA 0.248 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0812 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.1 2.625 2.5 3.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.76 -0.4 7.26 0.4 ;
      RECT 6.42 -0.4 6.76 0.95 ;
      RECT 5.32 -0.4 6.42 0.4 ;
      RECT 4.98 -0.4 5.32 1.115 ;
      RECT 0.52 -0.4 4.98 0.4 ;
      RECT 0.18 -0.4 0.52 1.465 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.355 4.64 7.26 5.44 ;
      RECT 5.965 4.465 6.355 5.44 ;
      RECT 4.445 4.64 5.965 5.44 ;
      RECT 4.105 4.465 4.445 5.44 ;
      RECT 2.84 4.64 4.105 5.44 ;
      RECT 2.5 4.465 2.84 5.44 ;
      RECT 1.3 4.64 2.5 5.44 ;
      RECT 0.91 4.465 1.3 5.44 ;
      RECT 0 4.64 0.91 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.47 2.13 5.715 2.47 ;
      RECT 5.24 1.38 5.47 3.195 ;
      RECT 4.455 1.38 5.24 1.61 ;
      RECT 4.74 2.965 5.24 3.195 ;
      RECT 4.51 2.965 4.74 4.195 ;
      RECT 3.625 3.965 4.51 4.195 ;
      RECT 4.225 1.065 4.455 1.61 ;
      RECT 2.92 1.065 4.225 1.295 ;
      RECT 3.285 3.965 3.625 4.365 ;
      RECT 2.08 3.965 3.285 4.195 ;
      RECT 2.58 1.01 2.92 1.35 ;
      RECT 1.74 3.965 2.08 4.365 ;
  END
END AND4X4

MACRO NAND2X0_HVT
  CLASS CORE ;
  FOREIGN NAND2X0_HVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ NAND2X0_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4335 ;
  ANTENNAPARTIALMETALAREA 0.7995 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8372 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.775 2.94 3.82 3.22 ;
      RECT 3.71 1.505 3.775 3.22 ;
      RECT 3.545 0.835 3.71 4.05 ;
      RECT 3.48 0.835 3.545 1.735 ;
      RECT 3.48 2.72 3.545 4.05 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2618 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2137 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.5 2.2 2.64 2.545 ;
      RECT 2.195 1.845 2.5 2.545 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2162 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2402 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.72 2.44 1.95 3.195 ;
      RECT 1.535 2.965 1.72 3.195 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2243 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.005 2.255 1.29 2.715 ;
      RECT 0.8 2.255 1.005 2.71 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2826 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1554 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.67 0.565 2.335 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.935 -0.4 3.96 0.4 ;
      RECT 2.595 -0.4 2.935 0.575 ;
      RECT 0 -0.4 2.595 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.015 4.64 3.96 5.44 ;
      RECT 2.605 4.405 3.015 5.44 ;
      RECT 1.85 4.64 2.605 5.44 ;
      RECT 1.51 4.465 1.85 5.44 ;
      RECT 0.57 4.64 1.51 5.44 ;
      RECT 0.175 4.465 0.57 5.44 ;
      RECT 0 4.64 0.175 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.2 1.985 3.31 2.335 ;
      RECT 2.97 0.885 3.2 3.735 ;
      RECT 0.56 0.885 2.97 1.115 ;
      RECT 0.75 3.505 2.97 3.735 ;
      RECT 0.275 0.885 0.56 1.44 ;
      RECT 0.22 1.05 0.275 1.44 ;
  END
END NAND2X0_HVT

MACRO AND4X1
  CLASS CORE ;
  FOREIGN AND4X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ NAND2X0_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7294 ;
  ANTENNAPARTIALMETALAREA 0.7751 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4821 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.76 3.195 3.82 3.8 ;
      RECT 3.53 1.025 3.76 3.8 ;
      RECT 3.42 1.025 3.53 1.365 ;
      RECT 3.44 3.195 3.53 3.8 ;
      RECT 3.42 3.36 3.44 3.8 ;
     END
  END Y

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2886 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1395 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.53 2.405 3.085 2.925 ;
     END
  END D

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2343 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0335 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.41 2.38 1.84 2.925 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.3382 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.63 1.675 1.18 2.29 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1368 ;
  ANTENNAPARTIALMETALAREA 0.2632 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1289 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.585 0.53 3.26 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3 -0.4 3.96 0.4 ;
      RECT 2.66 -0.4 3 0.575 ;
      RECT 0 -0.4 2.66 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.1 4.64 3.96 5.44 ;
      RECT 0.93 4.465 3.1 5.44 ;
      RECT 0 4.64 0.93 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 3.16 1.685 3.27 2.025 ;
      RECT 2.93 0.935 3.16 2.025 ;
      RECT 0.52 0.935 2.93 1.165 ;
      RECT 2.3 1.74 2.93 1.97 ;
      RECT 2.26 1.74 2.3 3.46 ;
      RECT 2.07 1.74 2.26 3.725 ;
      RECT 1.92 3.155 2.07 3.725 ;
      RECT 0.52 3.495 1.92 3.725 ;
      RECT 0.18 0.935 0.52 1.275 ;
  END
END AND4X1

MACRO AOI211XL
  CLASS CORE ;
  FOREIGN AOI211XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.9436 ;
  ANTENNAPARTIALMETALAREA 0.8429 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1287 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.93 1.15 3.16 3.195 ;
      RECT 1.46 1.15 2.93 1.38 ;
      RECT 2.78 2.965 2.93 3.195 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2337 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.51 2.33 2.125 2.71 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.252 ;
  ANTENNAPARTIALMETALAREA 0.2523 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.325 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.47 1.82 2.7 2.485 ;
      RECT 2.115 1.82 2.47 2.1 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.2679 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1501 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.955 0.52 2.66 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2772 ;
  ANTENNAPARTIALMETALAREA 0.261 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0918 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.795 1.65 1.375 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.46 -0.4 3.3 0.4 ;
      RECT 2.12 -0.4 2.46 0.575 ;
      RECT 0.52 -0.4 2.12 0.4 ;
      RECT 0.18 -0.4 0.52 1.24 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.08 4.64 3.3 5.44 ;
      RECT 0.74 4.465 1.08 5.44 ;
      RECT 0 4.64 0.74 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.18 2.955 1.84 3.185 ;
  END
END AOI211XL

MACRO AOI211X4
  CLASS CORE ;
  FOREIGN AOI211X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI211XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4374 ;
  ANTENNAPARTIALMETALAREA 0.8455 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1164 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.14 0.76 5.325 1.585 ;
      RECT 5.14 2.74 5.195 3.08 ;
      RECT 5.095 0.76 5.14 3.08 ;
      RECT 4.855 1.26 5.095 3.08 ;
      RECT 4.76 1.26 4.855 2.66 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.2524 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.305 2.38 2.07 2.71 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2268 ;
  ANTENNAPARTIALMETALAREA 0.3059 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2561 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.78 2.415 3.16 3.22 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.2282 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.215 1.285 0.495 2.1 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2484 ;
  ANTENNAPARTIALMETALAREA 0.208 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 1.775 1.44 2.1 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.1 -0.4 6.6 0.4 ;
      RECT 5.76 -0.4 6.1 1.42 ;
      RECT 4.66 -0.4 5.76 0.4 ;
      RECT 4.32 -0.4 4.66 0.895 ;
      RECT 2.34 -0.4 4.32 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 0.52 -0.4 2 0.4 ;
      RECT 0.18 -0.4 0.52 0.895 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.835 4.64 6.6 5.44 ;
      RECT 5.495 4.01 5.835 5.44 ;
      RECT 4.555 4.64 5.495 5.44 ;
      RECT 4.215 3.815 4.555 5.44 ;
      RECT 1.085 4.64 4.215 5.44 ;
      RECT 0.745 4.465 1.085 5.44 ;
      RECT 0 4.64 0.745 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.6 2.18 5.83 3.58 ;
      RECT 4.315 3.35 5.6 3.58 ;
      RECT 4.085 1.135 4.315 3.58 ;
      RECT 3.885 1.135 4.085 1.365 ;
      RECT 3.835 3.055 4.085 3.58 ;
      RECT 3.655 0.88 3.885 1.365 ;
      RECT 3.295 1.735 3.85 1.965 ;
      RECT 3.495 3.055 3.835 3.875 ;
      RECT 3.065 1.13 3.295 1.965 ;
      RECT 2.53 3.465 3.13 3.695 ;
      RECT 1.5 1.13 3.065 1.36 ;
      RECT 2.53 1.735 3.065 1.965 ;
      RECT 2.3 1.735 2.53 3.695 ;
      RECT 0.18 3.235 1.85 3.465 ;
  END
END AOI211X4

MACRO AOI211X2
  CLASS CORE ;
  FOREIGN AOI211X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.94 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI211XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.72 ;
  ANTENNAPARTIALMETALAREA 2.2638 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.1813 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.46 1.045 5.69 3.195 ;
      RECT 5.25 1.045 5.46 1.275 ;
      RECT 4.37 2.965 5.46 3.195 ;
      RECT 4.91 0.935 5.25 1.275 ;
      RECT 3.64 0.99 4.91 1.22 ;
      RECT 4.085 2.965 4.37 3.39 ;
      RECT 4.03 3.05 4.085 3.39 ;
      RECT 2.83 0.935 3.64 1.275 ;
      RECT 2.78 0.935 2.83 1.22 ;
      RECT 0.53 0.99 2.78 1.22 ;
      RECT 0.19 0.935 0.53 1.275 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.9051 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.2082 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.995 1.535 5.225 2.265 ;
      RECT 4.76 1.535 4.995 1.845 ;
      RECT 3.36 1.535 4.76 1.765 ;
      RECT 3.13 1.535 3.36 2.635 ;
      RECT 2.855 2.31 3.13 2.635 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.276 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1554 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.79 2.31 4.48 2.71 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.2238 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0335 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.265 1.48 2.635 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7986 ;
  ANTENNAPARTIALMETALAREA 0.7494 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4821 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.23 2.075 2.285 2.61 ;
      RECT 2 1.675 2.23 2.61 ;
      RECT 0.77 1.675 2 1.905 ;
      RECT 1.945 2.27 2 2.61 ;
      RECT 0.445 1.62 0.77 1.96 ;
      RECT 0.43 1.62 0.445 2.075 ;
      RECT 0.215 1.675 0.43 2.075 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 4.485 -0.4 5.94 0.4 ;
      RECT 4.145 -0.4 4.485 0.575 ;
      RECT 1.85 -0.4 4.145 0.4 ;
      RECT 1.51 -0.4 1.85 0.575 ;
      RECT 0 -0.4 1.51 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.445 4.64 5.94 5.44 ;
      RECT 2.105 3.82 2.445 5.44 ;
      RECT 1.165 4.64 2.105 5.44 ;
      RECT 0.825 3.82 1.165 5.44 ;
      RECT 0 4.64 0.825 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.31 3.7 5.65 4.04 ;
      RECT 3.48 3.755 5.31 3.985 ;
      RECT 3.25 2.89 3.48 3.985 ;
      RECT 0.185 2.89 3.25 3.12 ;
  END
END AOI211X2

MACRO AOI211X1
  CLASS CORE ;
  FOREIGN AOI211X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AOI211XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.366 ;
  ANTENNAPARTIALMETALAREA 1.3846 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.8989 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.08 1.095 3.18 3.195 ;
      RECT 3.01 1.095 3.08 4.095 ;
      RECT 2.95 0.805 3.01 4.095 ;
      RECT 2.78 0.805 2.95 1.435 ;
      RECT 2.74 2.775 2.95 4.095 ;
      RECT 1.835 0.805 2.78 1.035 ;
      RECT 1.605 0.805 1.835 1.38 ;
      RECT 1.46 1.15 1.605 1.38 ;
     END
  END Y

  PIN C0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.2895 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1448 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.165 2.045 2.66 ;
     END
  END C0

  PIN B0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.36 ;
  ANTENNAPARTIALMETALAREA 0.3818 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0034 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.51 1.83 2.72 2.25 ;
      RECT 2.49 1.83 2.51 3.195 ;
      RECT 2.28 2.02 2.49 3.195 ;
      RECT 2.195 2.965 2.28 3.195 ;
     END
  END B0

  PIN A1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4029 ;
  ANTENNAPARTIALMETALAREA 0.2575 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 2.2 0.645 2.71 ;
     END
  END A1

  PIN A0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4029 ;
  ANTENNAPARTIALMETALAREA 0.2481 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2508 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.68 1.43 1.91 ;
      RECT 0.875 1.285 1.18 1.91 ;
     END
  END A0

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.345 -0.4 3.3 0.4 ;
      RECT 2.005 -0.4 2.345 0.575 ;
      RECT 0.52 -0.4 2.005 0.4 ;
      RECT 0.18 -0.4 0.52 1.155 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.16 4.64 3.3 5.44 ;
      RECT 0.82 3.755 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 0.18 3.115 1.8 3.345 ;
  END
END AOI211X1

MACRO AND3XL
  CLASS CORE ;
  FOREIGN AND3XL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5694 ;
  ANTENNAPARTIALMETALAREA 0.8998 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.869 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.15 3.495 3.16 4.24 ;
      RECT 2.92 1.15 3.15 4.24 ;
      RECT 2.78 1.15 2.92 1.49 ;
      RECT 2.74 3.495 2.92 4.24 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1512 ;
  ANTENNAPARTIALMETALAREA 0.2236 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.455 1.715 1.975 2.145 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1512 ;
  ANTENNAPARTIALMETALAREA 0.2298 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.63 2.845 1.135 3.3 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1512 ;
  ANTENNAPARTIALMETALAREA 0.2244 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.79 0.58 2.3 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.34 -0.4 3.3 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 0 -0.4 2 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.465 4.64 3.3 5.44 ;
      RECT 2.465 2.62 2.69 3.125 ;
      RECT 2.235 2.62 2.465 5.44 ;
      RECT 1.34 4.64 2.235 5.44 ;
      RECT 1.335 4.465 1.34 5.44 ;
      RECT 1.01 4.41 1.335 5.44 ;
      RECT 1 4.465 1.01 5.44 ;
      RECT 0 4.64 1 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.55 1.75 2.69 2.1 ;
      RECT 2.32 1.125 2.55 2.1 ;
      RECT 1.055 1.125 2.32 1.355 ;
      RECT 1.52 2.38 1.75 4.18 ;
      RECT 1.465 2.38 1.52 3.125 ;
      RECT 0.54 3.95 1.52 4.18 ;
      RECT 1.055 2.38 1.465 2.61 ;
      RECT 0.825 1.125 1.055 2.61 ;
      RECT 0.52 1.125 0.825 1.355 ;
      RECT 0.2 3.95 0.54 4.355 ;
      RECT 0.18 1.07 0.52 1.41 ;
  END
END AND3XL

MACRO AND3X4
  CLASS CORE ;
  FOREIGN AND3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND3XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3307 ;
  ANTENNAPARTIALMETALAREA 1.011 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.71 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.745 1.82 3.82 3.22 ;
      RECT 3.44 1.69 3.745 3.22 ;
      RECT 2.985 1.69 3.44 1.92 ;
      RECT 2.85 2.8 3.44 3.155 ;
      RECT 2.755 1.375 2.985 1.92 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4812 ;
  ANTENNAPARTIALMETALAREA 0.243 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2773 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.835 1.82 2.065 2.42 ;
      RECT 1.46 1.82 1.835 2.1 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4812 ;
  ANTENNAPARTIALMETALAREA 0.2123 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.35 1.485 2.66 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4812 ;
  ANTENNAPARTIALMETALAREA 0.2601 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.82 0.57 2.425 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.78 -0.4 3.96 0.4 ;
      RECT 3.44 -0.4 3.78 0.575 ;
      RECT 2.39 -0.4 3.44 0.4 ;
      RECT 2.05 -0.4 2.39 1.03 ;
      RECT 0 -0.4 2.05 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.78 4.64 3.96 5.44 ;
      RECT 3.44 3.855 3.78 5.44 ;
      RECT 2.46 4.64 3.44 5.44 ;
      RECT 2.12 3.75 2.46 5.44 ;
      RECT 1.16 4.64 2.12 5.44 ;
      RECT 0.82 3.75 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.525 2.295 3.065 2.525 ;
      RECT 2.295 1.33 2.525 3.37 ;
      RECT 1.605 1.33 2.295 1.56 ;
      RECT 0.18 3.14 2.295 3.37 ;
      RECT 1.375 1.135 1.605 1.56 ;
      RECT 0.535 1.135 1.375 1.365 ;
      RECT 0.195 1.08 0.535 1.42 ;
  END
END AND3X4

MACRO AND3X2
  CLASS CORE ;
  FOREIGN AND3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND3XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3616 ;
  ANTENNAPARTIALMETALAREA 0.7263 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1747 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.96 1.33 3.1 3.195 ;
      RECT 2.87 0.79 2.96 3.195 ;
      RECT 2.62 0.79 2.87 1.61 ;
      RECT 2.815 2.74 2.87 3.195 ;
      RECT 2.76 2.74 2.815 3.08 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2664 ;
  ANTENNAPARTIALMETALAREA 0.3389 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.6907 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.87 2.52 1.98 2.895 ;
      RECT 1.64 1.82 1.87 2.895 ;
      RECT 1.46 1.82 1.64 2.1 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2664 ;
  ANTENNAPARTIALMETALAREA 0.2366 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.025 2.37 1.255 2.895 ;
      RECT 0.8 2.38 1.025 2.895 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2664 ;
  ANTENNAPARTIALMETALAREA 0.3134 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 2.465 0.57 2.805 ;
      RECT 0.14 2.465 0.52 3.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.2 -0.4 3.3 0.4 ;
      RECT 1.86 -0.4 2.2 0.575 ;
      RECT 0 -0.4 1.86 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.34 4.64 3.3 5.44 ;
      RECT 2 4.41 2.34 5.44 ;
      RECT 0 4.64 2 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.475 2.05 2.64 2.45 ;
      RECT 2.39 2.05 2.475 3.48 ;
      RECT 2.245 1.36 2.39 3.48 ;
      RECT 2.16 1.36 2.245 2.28 ;
      RECT 1.12 3.25 2.245 3.48 ;
      RECT 0.52 1.36 2.16 1.59 ;
      RECT 0.89 3.25 1.12 4.235 ;
      RECT 0.52 4.005 0.89 4.235 ;
      RECT 0.18 1.25 0.52 1.59 ;
      RECT 0.175 4.005 0.52 4.405 ;
  END
END AND3X2

MACRO AND3X1
  CLASS CORE ;
  FOREIGN AND3X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND3XL ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7008 ;
  ANTENNAPARTIALMETALAREA 0.8638 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8213 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.92 1.15 3.15 4.155 ;
      RECT 2.69 1.15 2.92 1.49 ;
      RECT 2.78 3.48 2.92 4.155 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2236 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.455 1.715 1.975 2.145 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2298 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.675 2.845 1.18 3.3 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2244 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.14 1.79 0.58 2.3 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.34 -0.4 3.3 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 0 -0.4 2 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.545 4.64 3.3 5.44 ;
      RECT 2.545 2.755 2.69 3.095 ;
      RECT 2.315 2.755 2.545 5.44 ;
      RECT 1.32 4.64 2.315 5.44 ;
      RECT 1.315 4.465 1.32 5.44 ;
      RECT 0.99 4.41 1.315 5.44 ;
      RECT 0.98 4.465 0.99 5.44 ;
      RECT 0 4.64 0.98 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 2.435 1.75 2.69 2.115 ;
      RECT 2.205 1.19 2.435 2.115 ;
      RECT 1.055 1.19 2.205 1.42 ;
      RECT 1.695 2.38 1.75 3.125 ;
      RECT 1.465 2.38 1.695 4.18 ;
      RECT 1.055 2.38 1.465 2.61 ;
      RECT 0.52 3.95 1.465 4.18 ;
      RECT 0.825 1.19 1.055 2.61 ;
      RECT 0.52 1.19 0.825 1.42 ;
      RECT 0.18 1.08 0.52 1.42 ;
      RECT 0.18 3.95 0.52 4.36 ;
  END
END AND3X1

MACRO AND2X1_LVT
  CLASS CORE ;
  FOREIGN AND2X1_LVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.6492 ;
  ANTENNAPARTIALMETALAREA 0.5247 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6288 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.355 2.38 2.5 2.66 ;
      RECT 2.125 1.445 2.355 3.55 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2204 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.825 2.37 1.205 2.95 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1332 ;
  ANTENNAPARTIALMETALAREA 0.2054 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.15 1.82 0.565 2.315 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.79 -0.4 2.64 0.4 ;
      RECT 1.45 -0.4 1.79 0.575 ;
      RECT 0 -0.4 1.45 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.4 4.64 2.64 5.44 ;
      RECT 0.46 4.465 1.4 5.44 ;
      RECT 0 4.64 0.46 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.66 0.82 1.89 3.475 ;
      RECT 0.52 0.82 1.66 1.05 ;
      RECT 0.8 3.245 1.66 3.475 ;
      RECT 0.46 3.19 0.8 3.53 ;
      RECT 0.18 0.765 0.52 1.105 ;
  END
END AND2X1_LVT

MACRO AND2X4
  CLASS CORE ;
  FOREIGN AND2X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND2X1_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4513 ;
  ANTENNAPARTIALMETALAREA 1.241 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8425 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.155 1.82 3.16 3.22 ;
      RECT 2.875 1.39 3.155 3.35 ;
      RECT 2.78 1.37 2.875 3.35 ;
      RECT 2.17 1.37 2.78 1.82 ;
      RECT 2.125 3.01 2.78 3.35 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4644 ;
  ANTENNAPARTIALMETALAREA 0.4482 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0087 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.18 1.98 1.375 2.36 ;
      RECT 1.145 1.98 1.18 3.3 ;
      RECT 0.95 2.13 1.145 3.3 ;
      RECT 0.8 2.635 0.95 3.3 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4581 ;
  ANTENNAPARTIALMETALAREA 0.2869 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2031 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 2.025 0.53 2.41 ;
      RECT 0.14 2.025 0.52 2.77 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.11 -0.4 3.3 0.4 ;
      RECT 2.77 -0.4 3.11 1.085 ;
      RECT 1.76 -0.4 2.77 0.4 ;
      RECT 1.42 -0.4 1.76 0.575 ;
      RECT 0 -0.4 1.42 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 3.11 4.64 3.3 5.44 ;
      RECT 2.77 3.775 3.11 5.44 ;
      RECT 1.785 4.64 2.77 5.44 ;
      RECT 1.445 4.465 1.785 5.44 ;
      RECT 0.535 4.64 1.445 5.44 ;
      RECT 0.17 4.465 0.535 5.44 ;
      RECT 0 4.64 0.17 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.845 2.09 2.43 2.43 ;
      RECT 1.645 1.485 1.845 2.82 ;
      RECT 1.615 1.485 1.645 3.82 ;
      RECT 0.52 1.485 1.615 1.715 ;
      RECT 1.415 2.59 1.615 3.82 ;
      RECT 0.74 3.59 1.415 3.82 ;
      RECT 0.18 1.44 0.52 1.78 ;
  END
END AND2X4

MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND2X1_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3972 ;
  ANTENNAPARTIALMETALAREA 1.0689 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1658 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.42 0.955 2.465 3.22 ;
      RECT 2.235 0.82 2.42 4.21 ;
      RECT 2.195 0.82 2.235 1.845 ;
      RECT 2.08 2.89 2.235 4.21 ;
      RECT 2.08 0.82 2.195 1.64 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2376 ;
  ANTENNAPARTIALMETALAREA 0.238 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0441 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 3.5 1.36 3.925 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2376 ;
  ANTENNAPARTIALMETALAREA 0.2887 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2349 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 2.115 0.76 2.455 ;
      RECT 0.14 2.115 0.52 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.66 -0.4 2.64 0.4 ;
      RECT 1.32 -0.4 1.66 0.575 ;
      RECT 0 -0.4 1.32 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.57 4.64 2.64 5.44 ;
      RECT 0.18 4.465 0.57 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.225 2.15 1.965 2.495 ;
      RECT 0.995 1.46 1.225 3.095 ;
      RECT 0.52 1.46 0.995 1.69 ;
      RECT 0.815 2.745 0.995 3.095 ;
      RECT 0.18 1.35 0.52 1.69 ;
  END
END AND2X2

MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.64 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AND2X1_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.756 ;
  ANTENNAPARTIALMETALAREA 0.7642 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.3337 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.355 2.38 2.5 2.66 ;
      RECT 2.355 1.345 2.41 1.845 ;
      RECT 2.355 3.075 2.41 3.895 ;
      RECT 2.125 1.345 2.355 3.895 ;
      RECT 2.12 1.345 2.125 1.845 ;
      RECT 2.07 3.075 2.125 3.895 ;
      RECT 2.07 1.345 2.12 1.685 ;
     END
  END Y

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1224 ;
  ANTENNAPARTIALMETALAREA 0.2407 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0547 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 2.315 1.215 2.895 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1224 ;
  ANTENNAPARTIALMETALAREA 0.2054 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.15 1.82 0.565 2.315 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.79 -0.4 2.64 0.4 ;
      RECT 1.45 -0.4 1.79 0.575 ;
      RECT 0 -0.4 1.45 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.755 4.64 2.64 5.44 ;
      RECT 1.31 4.465 1.755 5.44 ;
      RECT 0.79 4.64 1.31 5.44 ;
      RECT 0.45 4.465 0.79 5.44 ;
      RECT 0 4.64 0.45 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 1.835 1.935 1.885 2.355 ;
      RECT 1.605 0.82 1.835 3.475 ;
      RECT 0.52 0.82 1.605 1.05 ;
      RECT 1.595 1.935 1.605 2.355 ;
      RECT 0.79 3.245 1.605 3.475 ;
      RECT 0.45 3.19 0.79 3.53 ;
      RECT 0.18 0.765 0.52 1.105 ;
  END
END AND2X1

MACRO ADDHXL
  CLASS CORE ;
  FOREIGN ADDHXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.0706 ;
  ANTENNAPARTIALMETALAREA 1.024 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9608 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.355 2.965 4.405 3.205 ;
      RECT 4.125 1.625 4.355 3.205 ;
      RECT 3.49 1.625 4.125 1.855 ;
      RECT 3.41 2.975 4.125 3.205 ;
      RECT 3.26 1.095 3.49 1.855 ;
      RECT 3.18 2.975 3.41 3.685 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.512 ;
  ANTENNAPARTIALMETALAREA 0.8119 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.9856 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.025 1.845 7.045 2.075 ;
      RECT 6.795 0.63 7.025 3.845 ;
      RECT 6.5 3.615 6.795 3.845 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.522 ;
  ANTENNAPARTIALMETALAREA 1.6044 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.2928 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.95 3.93 5.745 4.16 ;
      RECT 3.605 2.135 3.835 2.74 ;
      RECT 2.95 2.51 3.605 2.74 ;
      RECT 2.72 2.51 2.95 4.16 ;
      RECT 2.12 2.865 2.72 3.22 ;
      RECT 1.775 2.865 2.12 3.095 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3312 ;
  ANTENNAPARTIALMETALAREA 0.2604 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.18 2.31 5.8 2.73 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.36 -0.4 7.26 0.4 ;
      RECT 6.02 -0.4 6.36 0.97 ;
      RECT 5.065 -0.4 6.02 0.4 ;
      RECT 4.725 -0.4 5.065 0.575 ;
      RECT 1.28 -0.4 4.725 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.275 4.64 7.26 5.44 ;
      RECT 5.935 4.465 6.275 5.44 ;
      RECT 4.745 4.64 5.935 5.44 ;
      RECT 4.405 4.465 4.745 5.44 ;
      RECT 1.28 4.64 4.405 5.44 ;
      RECT 0.94 4.465 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.3 2.81 6.54 3.215 ;
      RECT 6.07 1.39 6.3 3.215 ;
      RECT 5.885 1.39 6.07 1.62 ;
      RECT 5.45 2.985 6.07 3.215 ;
      RECT 5.22 2.985 5.45 3.685 ;
      RECT 4.71 1.155 4.94 3.685 ;
      RECT 4.21 1.155 4.71 1.385 ;
      RECT 3.845 3.455 4.71 3.685 ;
      RECT 3.98 0.63 4.21 1.385 ;
      RECT 2.995 0.63 3.98 0.86 ;
      RECT 2.765 0.63 2.995 2.135 ;
      RECT 1.39 1.905 2.765 2.135 ;
      RECT 2.3 0.635 2.53 1.035 ;
      RECT 2.255 3.58 2.485 4.235 ;
      RECT 0.925 1.265 2.425 1.495 ;
      RECT 0.465 0.805 2.3 1.035 ;
      RECT 0.465 4.005 2.255 4.235 ;
      RECT 1.535 3.545 1.84 3.775 ;
      RECT 1.305 2.985 1.535 3.775 ;
      RECT 1.16 1.905 1.39 2.67 ;
      RECT 0.925 2.985 1.305 3.215 ;
      RECT 0.695 1.265 0.925 3.215 ;
      RECT 0.235 0.805 0.465 4.235 ;
  END
END ADDHXL

MACRO ADDHX4
  CLASS CORE ;
  FOREIGN ADDHX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 18.48 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 6.1304 ;
  ANTENNAPARTIALMETALAREA 3.2938 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 14.2888 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.34 0.665 10.65 1.005 ;
      RECT 8.135 0.665 10.34 0.895 ;
      RECT 5.725 2.985 10.245 3.215 ;
      RECT 7.905 0.665 8.135 1.645 ;
      RECT 7.705 1.26 7.905 1.645 ;
      RECT 5.8 1.415 7.705 1.645 ;
      RECT 5.725 1.26 5.8 2.66 ;
      RECT 5.495 1.26 5.725 3.215 ;
      RECT 5.42 1.26 5.495 2.66 ;
      RECT 4.78 2.985 5.495 3.215 ;
      RECT 5.22 1.315 5.42 1.7 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3188 ;
  ANTENNAPARTIALMETALAREA 0.9448 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7895 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.53 2.38 17.68 3.78 ;
      RECT 17.3 1.42 17.53 3.78 ;
      RECT 17.11 1.42 17.3 1.65 ;
      RECT 16.655 2.795 17.3 3.025 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 3.4386 ;
  ANTENNAPARTIALMETALAREA 0.9345 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5103 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.44 1.945 9.955 2.175 ;
      RECT 8.425 1.945 8.44 2.595 ;
      RECT 8.195 1.945 8.425 2.635 ;
      RECT 8.135 2.365 8.195 2.635 ;
      RECT 6.39 2.365 8.135 2.595 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 3.4914 ;
  ANTENNAPARTIALMETALAREA 0.8314 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.0757 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.4 2.05 15.505 2.28 ;
      RECT 12.17 1.845 12.4 2.28 ;
      RECT 12.095 1.845 12.17 2.075 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 18.09 -0.4 18.48 0.4 ;
      RECT 17.75 -0.4 18.09 0.96 ;
      RECT 16.81 -0.4 17.75 0.4 ;
      RECT 16.47 -0.4 16.81 0.96 ;
      RECT 15.465 -0.4 16.47 0.4 ;
      RECT 15.125 -0.4 15.465 0.95 ;
      RECT 14.185 -0.4 15.125 0.4 ;
      RECT 13.845 -0.4 14.185 0.95 ;
      RECT 12.905 -0.4 13.845 0.4 ;
      RECT 12.565 -0.4 12.905 0.895 ;
      RECT 4.68 -0.4 12.565 0.4 ;
      RECT 4.34 -0.4 4.68 0.575 ;
      RECT 3.12 -0.4 4.34 0.4 ;
      RECT 2.78 -0.4 3.12 0.575 ;
      RECT 1.8 -0.4 2.78 0.4 ;
      RECT 1.46 -0.4 1.8 0.96 ;
      RECT 0.52 -0.4 1.46 0.4 ;
      RECT 0.18 -0.4 0.52 0.95 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 17.745 4.64 18.48 5.44 ;
      RECT 17.295 4.465 17.745 5.44 ;
      RECT 16.335 4.64 17.295 5.44 ;
      RECT 15.995 4.09 16.335 5.44 ;
      RECT 15.03 4.64 15.995 5.44 ;
      RECT 14.69 4.09 15.03 5.44 ;
      RECT 13.75 4.64 14.69 5.44 ;
      RECT 13.41 4.09 13.75 5.44 ;
      RECT 12.425 4.64 13.41 5.44 ;
      RECT 12.085 4.465 12.425 5.44 ;
      RECT 10.865 4.64 12.085 5.44 ;
      RECT 10.525 4.465 10.865 5.44 ;
      RECT 4.48 4.64 10.525 5.44 ;
      RECT 4.14 4.465 4.48 5.44 ;
      RECT 3.12 4.64 4.14 5.44 ;
      RECT 2.78 4.465 3.12 5.44 ;
      RECT 1.8 4.64 2.78 5.44 ;
      RECT 1.46 4.09 1.8 5.44 ;
      RECT 0.52 4.64 1.46 5.44 ;
      RECT 0.18 4.09 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 16.16 2.095 16.755 2.325 ;
      RECT 15.93 2.095 16.16 2.765 ;
      RECT 13.49 1.49 16.105 1.72 ;
      RECT 11.64 2.535 15.93 2.765 ;
      RECT 12.3 3.005 15.675 3.235 ;
      RECT 13.205 1.36 13.49 1.72 ;
      RECT 12.23 1.36 13.205 1.59 ;
      RECT 12.07 3.005 12.3 3.68 ;
      RECT 12 0.715 12.23 1.59 ;
      RECT 10.705 3.45 12.07 3.68 ;
      RECT 11.11 0.715 12 0.945 ;
      RECT 11.57 2.535 11.64 3.125 ;
      RECT 11.34 1.39 11.57 3.125 ;
      RECT 11.285 2.895 11.34 3.125 ;
      RECT 10.88 0.715 11.11 1.645 ;
      RECT 10.705 1.415 10.88 1.645 ;
      RECT 10.475 1.415 10.705 4.215 ;
      RECT 8.445 1.415 10.475 1.645 ;
      RECT 8.02 3.985 10.475 4.215 ;
      RECT 7.79 3.68 8.02 4.215 ;
      RECT 5.385 3.68 7.79 3.91 ;
      RECT 5.16 0.665 7.425 0.895 ;
      RECT 4.94 4.145 7.04 4.375 ;
      RECT 5.155 3.535 5.385 3.91 ;
      RECT 4.93 0.665 5.16 1.04 ;
      RECT 2.905 3.535 5.155 3.765 ;
      RECT 3.745 1.515 4.975 1.745 ;
      RECT 4.71 4.005 4.94 4.375 ;
      RECT 2.875 0.81 4.93 1.04 ;
      RECT 2.44 4.005 4.71 4.235 ;
      RECT 3.515 1.515 3.745 3.08 ;
      RECT 2.68 2.18 2.905 3.765 ;
      RECT 2.645 0.81 2.875 1.645 ;
      RECT 2.675 2.07 2.68 3.765 ;
      RECT 0.93 2.07 2.675 2.41 ;
      RECT 0.695 1.415 2.645 1.645 ;
      RECT 2.21 2.795 2.44 4.235 ;
      RECT 0.695 2.795 2.21 3.025 ;
      RECT 0.465 1.415 0.695 3.025 ;
  END
END ADDHX4

MACRO ADDHX2
  CLASS CORE ;
  FOREIGN ADDHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.88 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.8488 ;
  ANTENNAPARTIALMETALAREA 1.9694 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.1355 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.715 1.285 5.945 1.645 ;
      RECT 4.24 2.83 5.86 3.17 ;
      RECT 3.515 1.34 5.715 1.57 ;
      RECT 3.745 2.885 4.24 3.17 ;
      RECT 3.265 2.885 3.745 3.195 ;
      RECT 3.32 1.285 3.515 1.57 ;
      RECT 3.265 1.285 3.32 1.625 ;
      RECT 3.035 1.285 3.265 3.195 ;
      RECT 2.98 1.285 3.035 1.625 ;
      RECT 3.015 2.81 3.035 3.195 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2792 ;
  ANTENNAPARTIALMETALAREA 0.6283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8355 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.08 1.36 11.505 1.7 ;
      RECT 11.005 1.36 11.08 1.845 ;
      RECT 11.015 2.63 11.07 3.08 ;
      RECT 11.005 2.63 11.015 3.195 ;
      RECT 10.775 1.47 11.005 3.195 ;
      RECT 10.73 2.63 10.775 3.08 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.7286 ;
  ANTENNAPARTIALMETALAREA 0.5714 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6924 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.145 1.84 5.485 2.18 ;
      RECT 5.065 1.84 5.145 2.125 ;
      RECT 4.835 1.845 5.065 2.125 ;
      RECT 4.1 1.895 4.835 2.125 ;
      RECT 3.87 1.895 4.1 2.6 ;
      RECT 3.76 2.26 3.87 2.6 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.7748 ;
  ANTENNAPARTIALMETALAREA 0.6088 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.279 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.365 1.905 9.375 2.245 ;
      RECT 8.135 1.845 8.365 2.245 ;
      RECT 7.625 1.905 8.135 2.245 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.785 -0.4 11.88 0.4 ;
      RECT 10.445 -0.4 10.785 0.95 ;
      RECT 9.525 -0.4 10.445 0.4 ;
      RECT 9.185 -0.4 9.525 0.985 ;
      RECT 8.245 -0.4 9.185 0.4 ;
      RECT 7.905 -0.4 8.245 0.985 ;
      RECT 1.84 -0.4 7.905 0.4 ;
      RECT 1.5 -0.4 1.84 0.575 ;
      RECT 0.52 -0.4 1.5 0.4 ;
      RECT 0.18 -0.4 0.52 0.965 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.43 4.64 11.88 5.44 ;
      RECT 10.09 4.09 10.43 5.44 ;
      RECT 9.09 4.64 10.09 5.44 ;
      RECT 8.75 4.09 9.09 5.44 ;
      RECT 7.81 4.64 8.75 5.44 ;
      RECT 7.47 4.145 7.81 5.44 ;
      RECT 6.56 4.64 7.47 5.44 ;
      RECT 6.22 4.41 6.56 5.44 ;
      RECT 1.84 4.64 6.22 5.44 ;
      RECT 1.5 4.465 1.84 5.44 ;
      RECT 0.52 4.64 1.5 5.44 ;
      RECT 0.18 4.145 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 10.245 2.16 10.355 2.5 ;
      RECT 10.015 2.16 10.245 2.765 ;
      RECT 9.825 1.315 10.165 1.655 ;
      RECT 7.12 2.535 10.015 2.765 ;
      RECT 7.41 1.36 9.825 1.59 ;
      RECT 8.34 2.995 9.73 3.335 ;
      RECT 8.11 2.995 8.34 3.765 ;
      RECT 6.405 3.535 8.11 3.765 ;
      RECT 7.18 0.665 7.41 1.59 ;
      RECT 6.405 0.665 7.18 0.895 ;
      RECT 6.87 2.535 7.12 3.2 ;
      RECT 6.78 1.215 6.87 3.2 ;
      RECT 6.64 1.215 6.78 2.765 ;
      RECT 6.175 0.665 6.405 3.765 ;
      RECT 5.02 0.665 6.175 0.895 ;
      RECT 5.71 3.535 6.175 3.765 ;
      RECT 5.48 3.535 5.71 4.3 ;
      RECT 5.22 4.07 5.48 4.3 ;
      RECT 4.88 4.07 5.22 4.41 ;
      RECT 2.365 4.18 4.88 4.41 ;
      RECT 2.3 0.665 3.96 0.895 ;
      RECT 2.945 3.715 3.94 3.945 ;
      RECT 2.715 3.54 2.945 3.945 ;
      RECT 2.505 1.27 2.735 3.08 ;
      RECT 1.44 3.54 2.715 3.77 ;
      RECT 2.26 1.27 2.505 1.5 ;
      RECT 2.26 2.74 2.505 3.08 ;
      RECT 2.135 4 2.365 4.41 ;
      RECT 2.07 0.665 2.3 1.04 ;
      RECT 0.98 4 2.135 4.23 ;
      RECT 1.44 0.81 2.07 1.04 ;
      RECT 1.21 0.81 1.44 3.77 ;
      RECT 0.82 1.365 1.21 1.705 ;
      RECT 0.82 2.74 1.21 3.08 ;
      RECT 0.75 3.57 0.98 4.23 ;
      RECT 0.58 2.12 0.92 2.46 ;
      RECT 0.495 3.57 0.75 3.8 ;
      RECT 0.495 2.23 0.58 2.46 ;
      RECT 0.265 2.23 0.495 3.8 ;
  END
END ADDHX2

MACRO ADDHX1
  CLASS CORE ;
  FOREIGN ADDHX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.92 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.8762 ;
  ANTENNAPARTIALMETALAREA 1.1041 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.6481 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.005 1.33 4.235 3.22 ;
      RECT 3.59 1.33 4.005 1.56 ;
      RECT 3.245 2.84 4.005 3.22 ;
      RECT 3.36 1.21 3.59 1.56 ;
      RECT 3.015 2.84 3.245 3.73 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8148 ;
  ANTENNAPARTIALMETALAREA 0.752 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.71 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.61 1.845 7.705 2.075 ;
      RECT 7.4 1.38 7.61 2.075 ;
      RECT 7.38 1.38 7.4 3.115 ;
      RECT 7.17 1.845 7.38 3.115 ;
      RECT 7.025 2.885 7.17 3.115 ;
      RECT 6.795 2.885 7.025 3.97 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.846 ;
  ANTENNAPARTIALMETALAREA 2.1553 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.8103 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.835 2.52 6.065 3.445 ;
      RECT 5.16 3.215 5.835 3.445 ;
      RECT 4.93 3.215 5.16 4.235 ;
      RECT 2.785 4.005 4.93 4.235 ;
      RECT 3.545 1.8 3.775 2.52 ;
      RECT 2.785 2.29 3.545 2.52 ;
      RECT 2.555 2.29 2.785 4.235 ;
      RECT 2.195 2.29 2.555 2.66 ;
      RECT 2.115 2.29 2.195 2.575 ;
      RECT 1.775 2.235 2.115 2.575 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.846 ;
  ANTENNAPARTIALMETALAREA 0.2562 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0918 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.465 1.82 5.075 2.24 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.15 -0.4 7.92 0.4 ;
      RECT 6.92 -0.4 7.15 1.355 ;
      RECT 5.125 -0.4 6.92 0.4 ;
      RECT 6.815 1.125 6.92 1.355 ;
      RECT 6.585 1.125 6.815 1.72 ;
      RECT 4.785 -0.4 5.125 0.575 ;
      RECT 1.36 -0.4 4.785 0.4 ;
      RECT 1.02 -0.4 1.36 0.575 ;
      RECT 0 -0.4 1.02 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.48 4.64 7.92 5.44 ;
      RECT 6.14 4.465 6.48 5.44 ;
      RECT 4.78 4.64 6.14 5.44 ;
      RECT 4.44 4.465 4.78 5.44 ;
      RECT 1.28 4.64 4.44 5.44 ;
      RECT 0.94 4.465 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.525 1.98 6.84 2.32 ;
      RECT 6.35 0.665 6.69 0.895 ;
      RECT 6.35 1.98 6.525 3.905 ;
      RECT 6.295 0.665 6.35 3.905 ;
      RECT 6.12 0.665 6.295 2.21 ;
      RECT 5.625 3.675 6.295 3.905 ;
      RECT 5.6 1.21 5.885 1.55 ;
      RECT 5.395 3.675 5.625 4.04 ;
      RECT 5.545 1.21 5.6 2.985 ;
      RECT 5.37 1.265 5.545 2.985 ;
      RECT 4.7 1.265 5.37 1.495 ;
      RECT 4.7 2.755 5.37 2.985 ;
      RECT 4.47 0.805 4.7 1.495 ;
      RECT 4.47 2.755 4.7 3.775 ;
      RECT 4.365 0.805 4.47 1.035 ;
      RECT 3.68 3.545 4.47 3.775 ;
      RECT 4.025 0.675 4.365 1.035 ;
      RECT 3.13 0.675 4.025 0.905 ;
      RECT 2.9 0.675 3.13 1.955 ;
      RECT 1.385 1.725 2.9 1.955 ;
      RECT 2.44 0.63 2.67 1.035 ;
      RECT 0.925 1.265 2.55 1.495 ;
      RECT 0.465 0.805 2.44 1.035 ;
      RECT 2.095 4.005 2.325 4.405 ;
      RECT 0.465 4.005 2.095 4.235 ;
      RECT 1.5 3.18 1.84 3.52 ;
      RECT 0.925 3.18 1.5 3.41 ;
      RECT 1.155 1.725 1.385 2.56 ;
      RECT 0.695 1.265 0.925 3.41 ;
      RECT 0.235 0.76 0.465 4.235 ;
  END
END ADDHX1

MACRO ADDFXL
  CLASS CORE ;
  FOREIGN ADDFXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.7191 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0157 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.57 1.285 13.645 1.515 ;
      RECT 13.46 1.285 13.57 1.845 ;
      RECT 13.46 2.635 13.57 3.605 ;
      RECT 13.23 1.285 13.46 3.605 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.732 ;
  ANTENNAPARTIALMETALAREA 0.5743 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6235 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.005 2.38 12.325 2.66 ;
      RECT 11.985 1.43 12.005 2.66 ;
      RECT 11.755 1.43 11.985 3.135 ;
      RECT 11.665 1.43 11.755 1.77 ;
      RECT 11.645 2.795 11.755 3.135 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3816 ;
  ANTENNAPARTIALMETALAREA 0.5213 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4221 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.22 1.82 9.485 2.05 ;
      RECT 8.99 1.82 9.22 3.22 ;
      RECT 8.6 2.865 8.99 3.22 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5424 ;
  ANTENNAPARTIALMETALAREA 0.2214 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.04 0.76 2.38 ;
      RECT 0.42 2.04 0.445 2.635 ;
      RECT 0.215 2.15 0.42 2.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.54 ;
  ANTENNAPARTIALMETALAREA 0.3196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.895 2.35 4.835 2.69 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.77 -0.4 13.86 0.4 ;
      RECT 12.43 -0.4 12.77 1.615 ;
      RECT 10.08 -0.4 12.43 0.4 ;
      RECT 9.74 -0.4 10.08 0.575 ;
      RECT 4.725 -0.4 9.74 0.4 ;
      RECT 4.385 -0.4 4.725 0.9 ;
      RECT 1.285 -0.4 4.385 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.775 4.64 13.86 5.44 ;
      RECT 12.435 3.93 12.775 5.44 ;
      RECT 8.935 4.64 12.435 5.44 ;
      RECT 8.595 4.465 8.935 5.44 ;
      RECT 1.2 4.64 8.595 5.44 ;
      RECT 0.86 4.465 1.2 5.44 ;
      RECT 0 4.64 0.86 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.635 2.015 12.865 3.595 ;
      RECT 11.645 3.365 12.635 3.595 ;
      RECT 11.415 3.365 11.645 3.945 ;
      RECT 9.395 4.18 11.455 4.41 ;
      RECT 10.455 3.715 11.415 3.945 ;
      RECT 11.14 0.63 11.295 0.86 ;
      RECT 11.14 3.12 11.175 3.46 ;
      RECT 10.91 0.63 11.14 3.46 ;
      RECT 10.9 0.63 10.91 1.04 ;
      RECT 10.835 3.12 10.91 3.46 ;
      RECT 9.495 0.81 10.9 1.04 ;
      RECT 10.455 1.345 10.68 1.77 ;
      RECT 10.45 1.345 10.455 3.945 ;
      RECT 10.225 1.54 10.45 3.945 ;
      RECT 10.115 3.215 10.225 3.555 ;
      RECT 9.73 1.27 9.96 2.875 ;
      RECT 9.035 1.27 9.73 1.5 ;
      RECT 9.68 2.645 9.73 2.875 ;
      RECT 9.45 2.645 9.68 3.555 ;
      RECT 9.265 0.63 9.495 1.04 ;
      RECT 9.165 4.005 9.395 4.41 ;
      RECT 5.88 0.63 9.265 0.86 ;
      RECT 7.855 4.005 9.165 4.235 ;
      RECT 8.805 1.09 9.035 1.5 ;
      RECT 6.67 1.09 8.805 1.32 ;
      RECT 8.57 2.195 8.76 2.535 ;
      RECT 8.34 1.585 8.57 2.535 ;
      RECT 8.315 2.305 8.34 2.535 ;
      RECT 8.085 2.305 8.315 3.77 ;
      RECT 7.85 3.58 7.855 4.235 ;
      RECT 7.625 1.585 7.85 4.235 ;
      RECT 7.62 1.585 7.625 3.81 ;
      RECT 7.175 3.58 7.62 3.81 ;
      RECT 7.16 1.79 7.39 3.35 ;
      RECT 7.13 1.79 7.16 2.02 ;
      RECT 6.795 3.12 7.16 3.35 ;
      RECT 6.9 1.585 7.13 2.02 ;
      RECT 6.67 2.36 6.93 2.7 ;
      RECT 6.685 3.12 6.795 3.78 ;
      RECT 6.565 3.12 6.685 4.41 ;
      RECT 6.44 1.09 6.67 2.89 ;
      RECT 6.455 3.44 6.565 4.41 ;
      RECT 5.255 4.055 6.455 4.41 ;
      RECT 6.175 2.655 6.44 2.89 ;
      RECT 5.3 2.07 6.21 2.42 ;
      RECT 6.075 2.655 6.175 3.425 ;
      RECT 5.945 2.655 6.075 3.48 ;
      RECT 5.765 3.14 5.945 3.48 ;
      RECT 5.65 0.63 5.88 1.75 ;
      RECT 5.735 3.14 5.765 3.825 ;
      RECT 5.535 3.195 5.735 3.825 ;
      RECT 5.54 1.135 5.65 1.75 ;
      RECT 4.155 1.135 5.54 1.365 ;
      RECT 3.44 3.595 5.535 3.825 ;
      RECT 5.07 1.635 5.3 3.365 ;
      RECT 1.66 4.18 5.255 4.41 ;
      RECT 3.695 1.635 5.07 1.865 ;
      RECT 3.9 3.135 5.07 3.365 ;
      RECT 3.925 0.875 4.155 1.365 ;
      RECT 2.45 0.875 3.925 1.105 ;
      RECT 3.67 2.98 3.9 3.365 ;
      RECT 3.465 1.44 3.695 1.865 ;
      RECT 3.21 3.03 3.44 3.825 ;
      RECT 3.18 3.03 3.21 3.26 ;
      RECT 2.95 2.075 3.18 3.26 ;
      RECT 2.75 3.495 2.98 3.95 ;
      RECT 2.91 2.075 2.95 2.305 ;
      RECT 2.68 1.42 2.91 2.305 ;
      RECT 2.125 3.495 2.75 3.725 ;
      RECT 2.45 2.535 2.62 3.265 ;
      RECT 2.39 0.875 2.45 3.265 ;
      RECT 2.22 0.875 2.39 2.765 ;
      RECT 1.99 3.05 2.125 3.725 ;
      RECT 1.895 1.395 1.99 3.725 ;
      RECT 1.76 1.395 1.895 3.28 ;
      RECT 1.505 2.94 1.76 3.28 ;
      RECT 1.43 3.655 1.66 4.41 ;
      RECT 1.38 2.04 1.49 2.38 ;
      RECT 1.235 3.655 1.43 3.885 ;
      RECT 1.235 1.395 1.38 2.38 ;
      RECT 1.15 1.395 1.235 3.885 ;
      RECT 0.52 1.395 1.15 1.625 ;
      RECT 1.005 2.095 1.15 3.885 ;
      RECT 0.18 2.89 1.005 3.23 ;
      RECT 0.18 0.815 0.52 1.625 ;
  END
END ADDFXL

MACRO ADDFX4
  CLASS CORE ;
  FOREIGN ADDFX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.18 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3036 ;
  ANTENNAPARTIALMETALAREA 0.9635 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.5652 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.72 1.395 13.935 3.155 ;
      RECT 13.595 1.395 13.72 3.22 ;
      RECT 13.34 1.82 13.595 3.22 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3036 ;
  ANTENNAPARTIALMETALAREA 1.0169 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6076 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.4 1.395 12.655 3.155 ;
      RECT 12.315 1.395 12.4 3.22 ;
      RECT 12.02 1.82 12.315 3.22 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3816 ;
  ANTENNAPARTIALMETALAREA 0.5213 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4221 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.22 1.82 9.485 2.05 ;
      RECT 8.99 1.82 9.22 3.22 ;
      RECT 8.6 2.865 8.99 3.22 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5424 ;
  ANTENNAPARTIALMETALAREA 0.2214 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.04 0.76 2.38 ;
      RECT 0.42 2.04 0.445 2.635 ;
      RECT 0.215 2.15 0.42 2.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.54 ;
  ANTENNAPARTIALMETALAREA 0.3196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.895 2.35 4.835 2.69 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.575 -0.4 15.18 0.4 ;
      RECT 14.235 -0.4 14.575 1.005 ;
      RECT 13.295 -0.4 14.235 0.4 ;
      RECT 12.955 -0.4 13.295 1.005 ;
      RECT 12.015 -0.4 12.955 0.4 ;
      RECT 11.675 -0.4 12.015 1.005 ;
      RECT 10.08 -0.4 11.675 0.4 ;
      RECT 9.74 -0.4 10.08 0.575 ;
      RECT 4.725 -0.4 9.74 0.4 ;
      RECT 4.385 -0.4 4.725 0.905 ;
      RECT 1.285 -0.4 4.385 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.555 4.64 15.18 5.44 ;
      RECT 14.215 4.145 14.555 5.44 ;
      RECT 13.275 4.64 14.215 5.44 ;
      RECT 12.935 4.145 13.275 5.44 ;
      RECT 11.995 4.64 12.935 5.44 ;
      RECT 11.655 4.145 11.995 5.44 ;
      RECT 8.935 4.64 11.655 5.44 ;
      RECT 8.595 4.465 8.935 5.44 ;
      RECT 1.2 4.64 8.595 5.44 ;
      RECT 0.86 4.465 1.2 5.44 ;
      RECT 0 4.64 0.86 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 14.165 2.015 14.395 3.915 ;
      RECT 10.455 3.685 14.165 3.915 ;
      RECT 9.395 4.18 11.365 4.41 ;
      RECT 11.185 0.63 11.285 0.86 ;
      RECT 10.955 0.63 11.185 3.42 ;
      RECT 10.9 0.63 10.955 1.04 ;
      RECT 10.835 3.175 10.955 3.42 ;
      RECT 9.495 0.81 10.9 1.04 ;
      RECT 10.45 1.345 10.67 2.36 ;
      RECT 10.45 3.215 10.455 3.915 ;
      RECT 10.44 1.345 10.45 3.915 ;
      RECT 10.225 2.13 10.44 3.915 ;
      RECT 10.22 2.13 10.225 3.555 ;
      RECT 10.115 3.215 10.22 3.555 ;
      RECT 9.72 1.27 9.95 2.875 ;
      RECT 9.035 1.27 9.72 1.5 ;
      RECT 9.68 2.645 9.72 2.875 ;
      RECT 9.45 2.645 9.68 3.555 ;
      RECT 9.265 0.63 9.495 1.04 ;
      RECT 9.165 4.005 9.395 4.41 ;
      RECT 5.88 0.63 9.265 0.86 ;
      RECT 7.855 4.005 9.165 4.235 ;
      RECT 8.805 1.09 9.035 1.5 ;
      RECT 6.67 1.09 8.805 1.32 ;
      RECT 8.57 2.195 8.76 2.535 ;
      RECT 8.34 1.585 8.57 2.535 ;
      RECT 8.315 2.305 8.34 2.535 ;
      RECT 8.085 2.305 8.315 3.77 ;
      RECT 7.85 3.58 7.855 4.235 ;
      RECT 7.625 1.585 7.85 4.235 ;
      RECT 7.62 1.585 7.625 3.81 ;
      RECT 7.175 3.58 7.62 3.81 ;
      RECT 7.16 1.79 7.39 3.35 ;
      RECT 7.13 1.79 7.16 2.02 ;
      RECT 6.795 3.12 7.16 3.35 ;
      RECT 6.9 1.585 7.13 2.02 ;
      RECT 6.67 2.36 6.93 2.7 ;
      RECT 6.685 3.12 6.795 3.845 ;
      RECT 6.565 3.12 6.685 4.41 ;
      RECT 6.44 1.09 6.67 2.89 ;
      RECT 6.455 3.505 6.565 4.41 ;
      RECT 5.255 4.055 6.455 4.41 ;
      RECT 6.175 2.655 6.44 2.89 ;
      RECT 5.3 2.07 6.21 2.42 ;
      RECT 6.075 2.655 6.175 3.425 ;
      RECT 5.945 2.655 6.075 3.48 ;
      RECT 5.765 3.14 5.945 3.48 ;
      RECT 5.65 0.63 5.88 1.75 ;
      RECT 5.735 3.14 5.765 3.825 ;
      RECT 5.535 3.195 5.735 3.825 ;
      RECT 5.54 1.135 5.65 1.75 ;
      RECT 4.155 1.135 5.54 1.365 ;
      RECT 3.44 3.595 5.535 3.825 ;
      RECT 5.07 1.635 5.3 3.365 ;
      RECT 1.66 4.18 5.255 4.41 ;
      RECT 3.695 1.635 5.07 1.865 ;
      RECT 3.9 3.135 5.07 3.365 ;
      RECT 3.925 0.875 4.155 1.365 ;
      RECT 2.45 0.875 3.925 1.105 ;
      RECT 3.67 2.98 3.9 3.365 ;
      RECT 3.465 1.44 3.695 1.865 ;
      RECT 3.21 3.03 3.44 3.825 ;
      RECT 3.18 3.03 3.21 3.26 ;
      RECT 2.95 2.075 3.18 3.26 ;
      RECT 2.75 3.495 2.98 3.95 ;
      RECT 2.91 2.075 2.95 2.305 ;
      RECT 2.68 1.42 2.91 2.305 ;
      RECT 2.125 3.495 2.75 3.725 ;
      RECT 2.45 2.535 2.62 3.16 ;
      RECT 2.39 0.875 2.45 3.16 ;
      RECT 2.22 0.875 2.39 2.765 ;
      RECT 1.99 3.05 2.125 3.725 ;
      RECT 1.895 1.395 1.99 3.725 ;
      RECT 1.76 1.395 1.895 3.28 ;
      RECT 1.505 2.94 1.76 3.28 ;
      RECT 1.43 3.655 1.66 4.41 ;
      RECT 1.38 2.04 1.49 2.38 ;
      RECT 1.235 3.655 1.43 3.885 ;
      RECT 1.235 1.395 1.38 2.38 ;
      RECT 1.15 1.395 1.235 3.885 ;
      RECT 0.52 1.395 1.15 1.625 ;
      RECT 1.005 2.095 1.15 3.885 ;
      RECT 0.18 2.89 1.005 3.23 ;
      RECT 0.18 0.815 0.52 1.625 ;
  END
END ADDFX4

MACRO ADDFX2
  CLASS CORE ;
  FOREIGN ADDFX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2616 ;
  ANTENNAPARTIALMETALAREA 0.5805 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.7295 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.325 1.285 13.37 1.78 ;
      RECT 13.325 2.795 13.355 3.135 ;
      RECT 13.095 1.285 13.325 3.135 ;
      RECT 13.03 1.285 13.095 1.78 ;
      RECT 13.015 2.795 13.095 3.135 ;
      RECT 12.755 1.285 13.03 1.515 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2728 ;
  ANTENNAPARTIALMETALAREA 0.5738 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.65 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.76 1.43 12.005 1.77 ;
      RECT 11.76 2.795 11.985 3.135 ;
      RECT 11.53 1.43 11.76 3.135 ;
      RECT 11.435 2.405 11.53 2.635 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3816 ;
  ANTENNAPARTIALMETALAREA 0.5213 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4221 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.22 1.82 9.485 2.05 ;
      RECT 8.99 1.82 9.22 3.22 ;
      RECT 8.6 2.865 8.99 3.22 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5424 ;
  ANTENNAPARTIALMETALAREA 0.2214 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.04 0.76 2.38 ;
      RECT 0.42 2.04 0.445 2.635 ;
      RECT 0.215 2.15 0.42 2.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.54 ;
  ANTENNAPARTIALMETALAREA 0.3196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.895 2.35 4.835 2.69 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.69 -0.4 13.86 0.4 ;
      RECT 12.35 -0.4 12.69 0.575 ;
      RECT 10.08 -0.4 12.35 0.4 ;
      RECT 9.74 -0.4 10.08 0.575 ;
      RECT 4.725 -0.4 9.74 0.4 ;
      RECT 4.385 -0.4 4.725 0.9 ;
      RECT 1.285 -0.4 4.385 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.675 4.64 13.86 5.44 ;
      RECT 12.335 4.465 12.675 5.44 ;
      RECT 8.935 4.64 12.335 5.44 ;
      RECT 8.595 4.465 8.935 5.44 ;
      RECT 1.2 4.64 8.595 5.44 ;
      RECT 0.86 4.465 1.2 5.44 ;
      RECT 0 4.64 0.86 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.635 2.015 12.865 2.39 ;
      RECT 12.515 2.16 12.635 2.39 ;
      RECT 12.285 2.16 12.515 3.945 ;
      RECT 10.455 3.715 12.285 3.945 ;
      RECT 9.395 4.18 11.365 4.41 ;
      RECT 11.13 0.63 11.285 0.86 ;
      RECT 11.13 3.12 11.175 3.46 ;
      RECT 10.9 0.63 11.13 3.46 ;
      RECT 9.495 0.81 10.9 1.04 ;
      RECT 10.835 3.12 10.9 3.46 ;
      RECT 10.45 1.345 10.67 2.36 ;
      RECT 10.45 3.215 10.455 3.945 ;
      RECT 10.44 1.345 10.45 3.945 ;
      RECT 10.225 2.13 10.44 3.945 ;
      RECT 10.22 2.13 10.225 3.555 ;
      RECT 10.115 3.215 10.22 3.555 ;
      RECT 9.72 1.27 9.95 2.875 ;
      RECT 9.035 1.27 9.72 1.5 ;
      RECT 9.68 2.645 9.72 2.875 ;
      RECT 9.45 2.645 9.68 3.555 ;
      RECT 9.265 0.63 9.495 1.04 ;
      RECT 9.165 4.005 9.395 4.41 ;
      RECT 5.88 0.63 9.265 0.86 ;
      RECT 7.855 4.005 9.165 4.235 ;
      RECT 8.805 1.09 9.035 1.5 ;
      RECT 6.67 1.09 8.805 1.32 ;
      RECT 8.57 2.195 8.76 2.535 ;
      RECT 8.34 1.585 8.57 2.535 ;
      RECT 8.315 2.305 8.34 2.535 ;
      RECT 8.085 2.305 8.315 3.77 ;
      RECT 7.85 3.58 7.855 4.235 ;
      RECT 7.625 1.585 7.85 4.235 ;
      RECT 7.62 1.585 7.625 3.81 ;
      RECT 7.175 3.58 7.62 3.81 ;
      RECT 7.16 1.79 7.39 3.35 ;
      RECT 7.13 1.79 7.16 2.02 ;
      RECT 6.795 3.12 7.16 3.35 ;
      RECT 6.9 1.585 7.13 2.02 ;
      RECT 6.67 2.36 6.93 2.7 ;
      RECT 6.685 3.12 6.795 3.845 ;
      RECT 6.565 3.12 6.685 4.41 ;
      RECT 6.44 1.09 6.67 2.89 ;
      RECT 6.455 3.505 6.565 4.41 ;
      RECT 5.255 4.055 6.455 4.41 ;
      RECT 6.175 2.655 6.44 2.89 ;
      RECT 5.3 2.07 6.21 2.42 ;
      RECT 6.075 2.655 6.175 3.425 ;
      RECT 5.945 2.655 6.075 3.48 ;
      RECT 5.765 3.14 5.945 3.48 ;
      RECT 5.65 0.63 5.88 1.75 ;
      RECT 5.735 3.14 5.765 3.825 ;
      RECT 5.535 3.195 5.735 3.825 ;
      RECT 5.54 1.135 5.65 1.75 ;
      RECT 4.155 1.135 5.54 1.365 ;
      RECT 3.44 3.595 5.535 3.825 ;
      RECT 5.07 1.635 5.3 3.365 ;
      RECT 1.66 4.18 5.255 4.41 ;
      RECT 3.695 1.635 5.07 1.865 ;
      RECT 3.9 3.135 5.07 3.365 ;
      RECT 3.925 0.875 4.155 1.365 ;
      RECT 2.45 0.875 3.925 1.105 ;
      RECT 3.67 2.98 3.9 3.365 ;
      RECT 3.465 1.44 3.695 1.865 ;
      RECT 3.21 3.03 3.44 3.825 ;
      RECT 3.18 3.03 3.21 3.26 ;
      RECT 2.95 2.075 3.18 3.26 ;
      RECT 2.75 3.495 2.98 3.95 ;
      RECT 2.91 2.075 2.95 2.305 ;
      RECT 2.68 1.42 2.91 2.305 ;
      RECT 2.125 3.495 2.75 3.725 ;
      RECT 2.45 2.535 2.62 3.16 ;
      RECT 2.39 0.875 2.45 3.16 ;
      RECT 2.22 0.875 2.39 2.765 ;
      RECT 1.99 3.05 2.125 3.725 ;
      RECT 1.895 1.395 1.99 3.725 ;
      RECT 1.76 1.395 1.895 3.28 ;
      RECT 1.505 2.94 1.76 3.28 ;
      RECT 1.43 3.655 1.66 4.41 ;
      RECT 1.38 2.04 1.49 2.38 ;
      RECT 1.235 3.655 1.43 3.885 ;
      RECT 1.235 1.395 1.38 2.38 ;
      RECT 1.15 1.395 1.235 3.885 ;
      RECT 0.52 1.395 1.15 1.625 ;
      RECT 1.005 2.095 1.15 3.885 ;
      RECT 0.18 2.89 1.005 3.23 ;
      RECT 0.18 0.815 0.52 1.625 ;
  END
END ADDFX2

MACRO ADDFX1
  CLASS CORE ;
  FOREIGN ADDFX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.7191 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0157 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.57 1.285 13.645 1.515 ;
      RECT 13.46 1.285 13.57 1.845 ;
      RECT 13.46 2.635 13.57 3.605 ;
      RECT 13.23 1.285 13.46 3.605 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.732 ;
  ANTENNAPARTIALMETALAREA 0.5743 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6235 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.005 2.38 12.325 2.66 ;
      RECT 11.985 1.43 12.005 2.66 ;
      RECT 11.755 1.43 11.985 3.135 ;
      RECT 11.665 1.43 11.755 1.77 ;
      RECT 11.645 2.795 11.755 3.135 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3816 ;
  ANTENNAPARTIALMETALAREA 0.5213 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4221 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.22 1.82 9.485 2.05 ;
      RECT 8.99 1.82 9.22 3.22 ;
      RECT 8.6 2.865 8.99 3.22 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5424 ;
  ANTENNAPARTIALMETALAREA 0.2214 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.04 0.76 2.38 ;
      RECT 0.42 2.04 0.445 2.635 ;
      RECT 0.215 2.15 0.42 2.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.54 ;
  ANTENNAPARTIALMETALAREA 0.3196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.895 2.35 4.835 2.69 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.77 -0.4 13.86 0.4 ;
      RECT 12.43 -0.4 12.77 1.615 ;
      RECT 10.08 -0.4 12.43 0.4 ;
      RECT 9.74 -0.4 10.08 0.575 ;
      RECT 4.725 -0.4 9.74 0.4 ;
      RECT 4.385 -0.4 4.725 0.9 ;
      RECT 1.285 -0.4 4.385 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.775 4.64 13.86 5.44 ;
      RECT 12.435 3.93 12.775 5.44 ;
      RECT 8.935 4.64 12.435 5.44 ;
      RECT 8.595 4.465 8.935 5.44 ;
      RECT 1.2 4.64 8.595 5.44 ;
      RECT 0.86 4.465 1.2 5.44 ;
      RECT 0 4.64 0.86 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.635 2.015 12.865 3.595 ;
      RECT 11.645 3.365 12.635 3.595 ;
      RECT 11.415 3.365 11.645 3.945 ;
      RECT 9.395 4.18 11.455 4.41 ;
      RECT 10.455 3.715 11.415 3.945 ;
      RECT 11.14 0.63 11.295 0.86 ;
      RECT 11.14 3.12 11.175 3.46 ;
      RECT 10.91 0.63 11.14 3.46 ;
      RECT 10.9 0.63 10.91 1.04 ;
      RECT 10.835 3.12 10.91 3.46 ;
      RECT 9.495 0.81 10.9 1.04 ;
      RECT 10.455 1.345 10.68 1.77 ;
      RECT 10.45 1.345 10.455 3.945 ;
      RECT 10.225 1.54 10.45 3.945 ;
      RECT 10.115 3.215 10.225 3.555 ;
      RECT 9.73 1.27 9.96 2.875 ;
      RECT 9.035 1.27 9.73 1.5 ;
      RECT 9.68 2.645 9.73 2.875 ;
      RECT 9.45 2.645 9.68 3.555 ;
      RECT 9.265 0.63 9.495 1.04 ;
      RECT 9.165 4.005 9.395 4.41 ;
      RECT 5.88 0.63 9.265 0.86 ;
      RECT 7.855 4.005 9.165 4.235 ;
      RECT 8.805 1.09 9.035 1.5 ;
      RECT 6.67 1.09 8.805 1.32 ;
      RECT 8.57 2.195 8.76 2.535 ;
      RECT 8.34 1.585 8.57 2.535 ;
      RECT 8.315 2.305 8.34 2.535 ;
      RECT 8.085 2.305 8.315 3.77 ;
      RECT 7.85 3.58 7.855 4.235 ;
      RECT 7.625 1.585 7.85 4.235 ;
      RECT 7.62 1.585 7.625 3.81 ;
      RECT 7.175 3.58 7.62 3.81 ;
      RECT 7.16 1.79 7.39 3.35 ;
      RECT 7.13 1.79 7.16 2.02 ;
      RECT 6.795 3.12 7.16 3.35 ;
      RECT 6.9 1.585 7.13 2.02 ;
      RECT 6.67 2.36 6.93 2.7 ;
      RECT 6.685 3.12 6.795 3.78 ;
      RECT 6.565 3.12 6.685 4.41 ;
      RECT 6.44 1.09 6.67 2.89 ;
      RECT 6.455 3.44 6.565 4.41 ;
      RECT 5.255 4.055 6.455 4.41 ;
      RECT 6.175 2.655 6.44 2.89 ;
      RECT 5.3 2.07 6.21 2.42 ;
      RECT 6.075 2.655 6.175 3.425 ;
      RECT 5.945 2.655 6.075 3.48 ;
      RECT 5.765 3.14 5.945 3.48 ;
      RECT 5.65 0.63 5.88 1.75 ;
      RECT 5.735 3.14 5.765 3.825 ;
      RECT 5.535 3.195 5.735 3.825 ;
      RECT 5.54 1.135 5.65 1.75 ;
      RECT 4.155 1.135 5.54 1.365 ;
      RECT 3.44 3.595 5.535 3.825 ;
      RECT 5.07 1.635 5.3 3.365 ;
      RECT 1.66 4.18 5.255 4.41 ;
      RECT 3.695 1.635 5.07 1.865 ;
      RECT 3.9 3.135 5.07 3.365 ;
      RECT 3.925 0.875 4.155 1.365 ;
      RECT 2.45 0.875 3.925 1.105 ;
      RECT 3.67 2.98 3.9 3.365 ;
      RECT 3.465 1.44 3.695 1.865 ;
      RECT 3.21 3.03 3.44 3.825 ;
      RECT 3.18 3.03 3.21 3.26 ;
      RECT 2.95 2.075 3.18 3.26 ;
      RECT 2.75 3.495 2.98 3.95 ;
      RECT 2.91 2.075 2.95 2.305 ;
      RECT 2.68 1.42 2.91 2.305 ;
      RECT 2.125 3.495 2.75 3.725 ;
      RECT 2.45 2.535 2.62 3.265 ;
      RECT 2.39 0.875 2.45 3.265 ;
      RECT 2.22 0.875 2.39 2.765 ;
      RECT 1.99 3.05 2.125 3.725 ;
      RECT 1.895 1.395 1.99 3.725 ;
      RECT 1.76 1.395 1.895 3.28 ;
      RECT 1.505 2.94 1.76 3.28 ;
      RECT 1.43 3.655 1.66 4.41 ;
      RECT 1.38 2.04 1.49 2.38 ;
      RECT 1.235 3.655 1.43 3.885 ;
      RECT 1.235 1.395 1.38 2.38 ;
      RECT 1.15 1.395 1.235 3.885 ;
      RECT 0.52 1.395 1.15 1.625 ;
      RECT 1.005 2.095 1.15 3.885 ;
      RECT 0.18 2.89 1.005 3.23 ;
      RECT 0.18 0.815 0.52 1.625 ;
  END
END ADDFX1

MACRO ADDFHXL
  CLASS CORE ;
  FOREIGN ADDFHXL 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.52 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 0.6181 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.7401 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.23 1.285 14.34 2.1 ;
      RECT 14.23 3.08 14.34 3.42 ;
      RECT 14 1.285 14.23 3.42 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.5088 ;
  ANTENNAPARTIALMETALAREA 0.6817 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1429 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.725 1.285 12.865 1.625 ;
      RECT 12.725 3.08 12.78 3.42 ;
      RECT 12.495 1.285 12.725 3.42 ;
      RECT 12.44 2.94 12.495 3.42 ;
      RECT 12.09 2.94 12.44 3.22 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1296 ;
  ANTENNAPARTIALMETALAREA 0.2098 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9858 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.36 2.675 11.745 3.22 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6336 ;
  ANTENNAPARTIALMETALAREA 0.2381 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1925 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.49 2.805 6.54 3.145 ;
      RECT 6.385 2.66 6.49 3.145 ;
      RECT 6.155 2.405 6.385 3.145 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2592 ;
  ANTENNAPARTIALMETALAREA 0.2515 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.75 2.085 1.18 2.67 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.625 -0.4 14.52 0.4 ;
      RECT 13.285 -0.4 13.625 0.575 ;
      RECT 12.255 -0.4 13.285 0.4 ;
      RECT 11.915 -0.4 12.255 0.575 ;
      RECT 6.955 -0.4 11.915 0.4 ;
      RECT 6.615 -0.4 6.955 0.575 ;
      RECT 1.32 -0.4 6.615 0.4 ;
      RECT 0.98 -0.4 1.32 0.575 ;
      RECT 0 -0.4 0.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.56 4.64 14.52 5.44 ;
      RECT 13.22 4.465 13.56 5.44 ;
      RECT 10.94 4.64 13.22 5.44 ;
      RECT 10.6 4.465 10.94 5.44 ;
      RECT 6.16 4.64 10.6 5.44 ;
      RECT 5.82 4.465 6.16 5.44 ;
      RECT 1.24 4.64 5.82 5.44 ;
      RECT 0.9 3.76 1.24 5.44 ;
      RECT 0 4.64 0.9 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.42 2.4 13.76 2.74 ;
      RECT 13.24 2.51 13.42 2.74 ;
      RECT 13.01 2.51 13.24 4.23 ;
      RECT 11.68 0.81 13.085 1.04 ;
      RECT 9.66 4 13.01 4.23 ;
      RECT 11.82 1.355 12.16 1.695 ;
      RECT 10.92 3.45 11.915 3.68 ;
      RECT 11.22 1.465 11.82 1.695 ;
      RECT 11.45 0.63 11.68 1.04 ;
      RECT 8.94 0.63 11.45 0.86 ;
      RECT 10.99 1.09 11.22 2.425 ;
      RECT 9.4 1.09 10.99 1.32 ;
      RECT 10.92 2.195 10.99 2.425 ;
      RECT 10.69 2.195 10.92 3.68 ;
      RECT 10.46 1.55 10.76 1.78 ;
      RECT 10.23 1.55 10.46 3.675 ;
      RECT 10.04 3.335 10.23 3.675 ;
      RECT 9.86 1.55 9.995 1.78 ;
      RECT 9.66 1.55 9.86 2.76 ;
      RECT 9.63 1.55 9.66 4.23 ;
      RECT 9.43 2.53 9.63 4.23 ;
      RECT 9.32 3.545 9.43 3.885 ;
      RECT 9.17 1.09 9.4 1.78 ;
      RECT 8.885 1.55 9.17 1.78 ;
      RECT 8.71 0.63 8.94 1.32 ;
      RECT 8.655 1.55 8.885 3.885 ;
      RECT 8.42 1.09 8.71 1.32 ;
      RECT 7.96 0.63 8.475 0.86 ;
      RECT 8.19 1.09 8.42 3.83 ;
      RECT 8.12 3.6 8.19 3.83 ;
      RECT 7.78 3.6 8.12 3.94 ;
      RECT 7.73 0.63 7.96 3.13 ;
      RECT 6.385 0.805 7.73 1.035 ;
      RECT 7.64 2.755 7.73 3.13 ;
      RECT 7.41 1.265 7.5 1.605 ;
      RECT 7.18 1.265 7.41 3.62 ;
      RECT 5.815 3.39 7.18 3.62 ;
      RECT 6.72 1.325 6.95 2.34 ;
      RECT 5.92 1.325 6.72 1.555 ;
      RECT 6.155 0.63 6.385 1.035 ;
      RECT 4.43 0.63 6.155 0.86 ;
      RECT 5.69 1.09 5.92 1.555 ;
      RECT 5.585 2.175 5.815 3.62 ;
      RECT 4.89 1.09 5.69 1.32 ;
      RECT 5.35 1.6 5.46 1.94 ;
      RECT 5.12 1.6 5.35 4.41 ;
      RECT 2.19 4.18 5.12 4.41 ;
      RECT 4.81 1.09 4.89 1.885 ;
      RECT 4.66 1.09 4.81 3.95 ;
      RECT 4.58 1.655 4.66 3.95 ;
      RECT 2.965 3.72 4.58 3.95 ;
      RECT 4.35 0.63 4.43 1.42 ;
      RECT 4.2 0.63 4.35 3.465 ;
      RECT 4.12 1.04 4.2 3.465 ;
      RECT 3.71 1.09 3.765 1.43 ;
      RECT 3.63 0.63 3.71 1.43 ;
      RECT 3.63 3.125 3.685 3.465 ;
      RECT 3.4 0.63 3.63 3.465 ;
      RECT 1.81 0.63 3.4 0.86 ;
      RECT 3.345 3.125 3.4 3.465 ;
      RECT 2.91 1.09 3.045 1.43 ;
      RECT 2.91 3.18 2.965 3.95 ;
      RECT 2.735 1.09 2.91 3.95 ;
      RECT 2.68 1.09 2.735 3.52 ;
      RECT 2.625 3.18 2.68 3.52 ;
      RECT 2.19 1.09 2.27 3.475 ;
      RECT 2.04 1.09 2.19 4.41 ;
      RECT 1.96 3.1 2.04 4.41 ;
      RECT 1.58 0.63 1.81 1.035 ;
      RECT 1.715 2.345 1.78 2.715 ;
      RECT 1.485 1.555 1.715 3.165 ;
      RECT 0.52 0.805 1.58 1.035 ;
      RECT 0.87 1.555 1.485 1.785 ;
      RECT 0.87 2.935 1.485 3.165 ;
      RECT 0.64 1.31 0.87 1.785 ;
      RECT 0.64 2.935 0.87 3.3 ;
      RECT 0.41 0.665 0.52 1.035 ;
      RECT 0.41 3.76 0.52 4.1 ;
      RECT 0.18 0.665 0.41 4.1 ;
  END
END ADDFHXL

MACRO ADDFHX4
  CLASS CORE ;
  FOREIGN ADDFHX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 23.1 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3188 ;
  ANTENNAPARTIALMETALAREA 0.7714 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.7772 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.15 1.82 22.3 3.22 ;
      RECT 21.92 1.4 22.15 3.22 ;
      RECT 21.71 1.4 21.92 1.74 ;
      RECT 21.71 2.82 21.92 3.16 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3212 ;
  ANTENNAPARTIALMETALAREA 0.7145 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6394 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.83 1.82 20.98 3.22 ;
      RECT 20.6 1.455 20.83 3.22 ;
      RECT 20.43 1.455 20.6 1.685 ;
      RECT 20.425 2.82 20.6 3.16 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6048 ;
  ANTENNAPARTIALMETALAREA 0.256 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.995 2.38 19.66 2.765 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.3112 ;
  ANTENNAPARTIALMETALAREA 0.4789 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.9186 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.645 2.665 14.07 3.005 ;
      RECT 13.415 2.665 13.645 3.195 ;
      RECT 12.79 2.665 13.415 3.005 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9162 ;
  ANTENNAPARTIALMETALAREA 0.3016 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.725 1.82 1.245 2.4 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 22.69 -0.4 23.1 0.4 ;
      RECT 22.35 -0.4 22.69 1.04 ;
      RECT 21.41 -0.4 22.35 0.4 ;
      RECT 21.07 -0.4 21.41 1.04 ;
      RECT 20.05 -0.4 21.07 0.4 ;
      RECT 19.71 -0.4 20.05 0.575 ;
      RECT 13.58 -0.4 19.71 0.4 ;
      RECT 13.24 -0.4 13.58 0.575 ;
      RECT 3.27 -0.4 13.24 0.4 ;
      RECT 2.93 -0.4 3.27 0.575 ;
      RECT 1.25 -0.4 2.93 0.4 ;
      RECT 0.91 -0.4 1.25 0.575 ;
      RECT 0 -0.4 0.91 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 22.695 4.64 23.1 5.44 ;
      RECT 22.355 4.085 22.695 5.44 ;
      RECT 21.41 4.64 22.355 5.44 ;
      RECT 21.07 4.085 21.41 5.44 ;
      RECT 20.125 4.64 21.07 5.44 ;
      RECT 19.785 4.09 20.125 5.44 ;
      RECT 18.815 4.64 19.785 5.44 ;
      RECT 18.365 4.465 18.815 5.44 ;
      RECT 14.09 4.64 18.365 5.44 ;
      RECT 13.75 4.01 14.09 5.44 ;
      RECT 12.65 4.64 13.75 5.44 ;
      RECT 12.31 4.01 12.65 5.44 ;
      RECT 3.66 4.64 12.31 5.44 ;
      RECT 3.32 3.765 3.66 5.44 ;
      RECT 1.445 4.64 3.32 5.44 ;
      RECT 1.105 4 1.445 5.44 ;
      RECT 0 4.64 1.105 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 21.44 2.21 21.625 2.58 ;
      RECT 21.21 2.21 21.44 3.835 ;
      RECT 17.265 3.605 21.21 3.835 ;
      RECT 20.305 2.025 20.36 2.365 ;
      RECT 20.02 1.915 20.305 2.365 ;
      RECT 19.91 1.915 20.02 2.145 ;
      RECT 19.68 1.005 19.91 2.145 ;
      RECT 19.055 1.005 19.68 1.235 ;
      RECT 18.59 1.495 19.45 1.725 ;
      RECT 18.59 3.045 19.365 3.275 ;
      RECT 18.825 0.63 19.055 1.235 ;
      RECT 15.965 0.63 18.825 0.86 ;
      RECT 18.36 1.09 18.59 3.275 ;
      RECT 16.49 1.09 18.36 1.32 ;
      RECT 18.165 2.305 18.36 2.67 ;
      RECT 17.93 1.55 18.13 1.78 ;
      RECT 17.93 2.99 17.985 3.33 ;
      RECT 17.7 1.55 17.93 3.33 ;
      RECT 17.645 2.99 17.7 3.33 ;
      RECT 17.21 1.55 17.405 1.78 ;
      RECT 17.21 3.295 17.265 4.105 ;
      RECT 16.98 1.55 17.21 4.105 ;
      RECT 16.925 3.295 16.98 4.105 ;
      RECT 16.49 3.155 16.545 3.965 ;
      RECT 16.26 1.09 16.49 3.965 ;
      RECT 16.205 3.155 16.26 3.965 ;
      RECT 15.91 0.63 15.965 1.52 ;
      RECT 15.68 0.63 15.91 3.43 ;
      RECT 15.625 0.7 15.68 1.52 ;
      RECT 15.66 3.2 15.68 3.43 ;
      RECT 15.32 3.2 15.66 4.02 ;
      RECT 15.165 0.635 15.395 2.88 ;
      RECT 15.15 0.635 15.165 1.035 ;
      RECT 12.745 0.805 15.15 1.035 ;
      RECT 14.81 1.46 14.935 3.68 ;
      RECT 14.705 1.46 14.81 4.31 ;
      RECT 14.34 1.46 14.705 1.69 ;
      RECT 14.47 3.45 14.705 4.31 ;
      RECT 14.245 1.92 14.475 2.29 ;
      RECT 13.37 3.45 14.47 3.68 ;
      RECT 14 1.35 14.34 1.69 ;
      RECT 13.26 1.92 14.245 2.15 ;
      RECT 13.03 3.45 13.37 4.31 ;
      RECT 13.03 1.265 13.26 2.15 ;
      RECT 12.195 1.265 13.03 1.495 ;
      RECT 12.195 3.45 13.03 3.68 ;
      RECT 12.195 1.725 12.78 1.955 ;
      RECT 12.515 0.66 12.745 1.035 ;
      RECT 9.705 0.66 12.515 0.89 ;
      RECT 11.965 1.13 12.195 1.495 ;
      RECT 11.965 1.725 12.195 3.78 ;
      RECT 10.165 1.13 11.965 1.36 ;
      RECT 11.505 1.595 11.735 4.295 ;
      RECT 10.395 1.595 11.505 1.825 ;
      RECT 9.97 4.065 11.505 4.295 ;
      RECT 11.035 2.06 11.265 3.815 ;
      RECT 10.165 2.06 11.035 2.29 ;
      RECT 7.24 3.585 11.035 3.815 ;
      RECT 10.58 3.1 10.785 3.33 ;
      RECT 10.35 2.525 10.58 3.33 ;
      RECT 9.705 2.525 10.35 2.755 ;
      RECT 9.935 1.13 10.165 2.29 ;
      RECT 9.685 4.065 9.97 4.34 ;
      RECT 9.475 0.63 9.705 2.755 ;
      RECT 4.38 4.11 9.685 4.34 ;
      RECT 9.19 3.095 9.48 3.325 ;
      RECT 8.34 0.63 9.475 0.86 ;
      RECT 8.96 1.26 9.19 3.325 ;
      RECT 8.72 1.26 8.96 1.49 ;
      RECT 7.815 3.095 8.96 3.325 ;
      RECT 8.285 2.635 8.72 2.865 ;
      RECT 8.285 0.63 8.34 1.33 ;
      RECT 8.11 0.63 8.285 2.865 ;
      RECT 8.055 0.99 8.11 2.865 ;
      RECT 8 0.99 8.055 1.33 ;
      RECT 7.585 1.95 7.815 3.325 ;
      RECT 7.565 0.99 7.62 1.33 ;
      RECT 7.565 1.95 7.585 2.18 ;
      RECT 7.51 0.99 7.565 2.18 ;
      RECT 7.335 0.63 7.51 2.18 ;
      RECT 7.28 0.63 7.335 1.33 ;
      RECT 6.175 0.63 7.28 0.86 ;
      RECT 7.185 3.045 7.24 3.865 ;
      RECT 6.98 2.46 7.185 3.865 ;
      RECT 6.955 1.185 6.98 3.865 ;
      RECT 6.75 1.185 6.955 2.69 ;
      RECT 6.9 3.045 6.955 3.865 ;
      RECT 5.045 3.635 6.9 3.865 ;
      RECT 6.56 1.185 6.75 1.415 ;
      RECT 6.39 3.095 6.52 3.325 ;
      RECT 6.16 2.4 6.39 3.325 ;
      RECT 6.12 0.63 6.175 1.13 ;
      RECT 6.12 2.4 6.16 2.63 ;
      RECT 5.89 0.63 6.12 2.63 ;
      RECT 5.835 0.63 5.89 1.13 ;
      RECT 3.735 0.63 5.835 0.86 ;
      RECT 5.51 3.1 5.82 3.33 ;
      RECT 5.48 1.605 5.51 3.33 ;
      RECT 5.425 1.55 5.48 3.33 ;
      RECT 5.28 1.09 5.425 3.33 ;
      RECT 5.195 1.09 5.28 1.92 ;
      RECT 4.2 1.09 5.195 1.32 ;
      RECT 5.14 1.55 5.195 1.89 ;
      RECT 4.815 2.505 5.045 3.865 ;
      RECT 4.695 2.505 4.815 2.735 ;
      RECT 4.465 1.55 4.695 2.735 ;
      RECT 4.15 3.1 4.38 4.34 ;
      RECT 4.03 1.09 4.2 1.685 ;
      RECT 4.04 3.1 4.15 3.985 ;
      RECT 3.78 3.1 4.04 3.53 ;
      RECT 3.97 1.09 4.03 1.74 ;
      RECT 3.78 1.4 3.97 1.74 ;
      RECT 3.69 1.4 3.78 3.53 ;
      RECT 3.505 0.63 3.735 1.04 ;
      RECT 3.55 1.455 3.69 3.53 ;
      RECT 2.71 1.455 3.55 1.685 ;
      RECT 2.94 3.3 3.55 3.53 ;
      RECT 0.52 0.81 3.505 1.04 ;
      RECT 2.85 2.09 3.19 2.43 ;
      RECT 2.6 3.3 2.94 3.64 ;
      RECT 1.955 2.145 2.85 2.375 ;
      RECT 2.37 1.4 2.71 1.74 ;
      RECT 1.965 4.055 2.4 4.285 ;
      RECT 1.955 1.46 2.01 1.8 ;
      RECT 1.735 3.45 1.965 4.285 ;
      RECT 1.785 1.46 1.955 2.375 ;
      RECT 1.785 2.74 1.84 3.08 ;
      RECT 1.725 1.46 1.785 3.08 ;
      RECT 0.52 3.45 1.735 3.68 ;
      RECT 1.67 1.46 1.725 1.8 ;
      RECT 1.555 2.145 1.725 3.08 ;
      RECT 1.5 2.74 1.555 3.08 ;
      RECT 0.465 0.81 0.52 1.63 ;
      RECT 0.465 2.83 0.52 4.25 ;
      RECT 0.29 0.81 0.465 4.25 ;
      RECT 0.235 1.29 0.29 4.25 ;
      RECT 0.18 1.29 0.235 1.63 ;
      RECT 0.18 2.83 0.235 4.25 ;
  END
END ADDFHX4

MACRO ADDFHX2
  CLASS CORE ;
  FOREIGN ADDFHX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.44 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4208 ;
  ANTENNAPARTIALMETALAREA 1.0283 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8425 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.05 0.92 22.23 2.075 ;
      RECT 22.05 2.635 22.105 4.025 ;
      RECT 21.89 0.92 22.05 4.025 ;
      RECT 21.82 1.5 21.89 4.025 ;
      RECT 21.765 2.745 21.82 4.025 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.0816 ;
  ANTENNAPARTIALMETALAREA 0.5978 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9256 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.79 1.39 20.97 1.73 ;
      RECT 20.63 1.39 20.79 3.195 ;
      RECT 20.56 1.445 20.63 3.195 ;
      RECT 20.015 2.965 20.56 3.195 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6048 ;
  ANTENNAPARTIALMETALAREA 0.2859 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1607 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.995 2.295 19.66 2.725 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.3112 ;
  ANTENNAPARTIALMETALAREA 0.4789 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.9186 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.645 2.665 14.07 3.005 ;
      RECT 13.415 2.665 13.645 3.195 ;
      RECT 12.79 2.665 13.415 3.005 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9162 ;
  ANTENNAPARTIALMETALAREA 0.3016 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.166 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.725 1.82 1.245 2.4 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 21.51 -0.4 22.44 0.4 ;
      RECT 21.17 -0.4 21.51 0.95 ;
      RECT 20.21 -0.4 21.17 0.4 ;
      RECT 19.87 -0.4 20.21 0.575 ;
      RECT 13.58 -0.4 19.87 0.4 ;
      RECT 13.24 -0.4 13.58 0.575 ;
      RECT 3.35 -0.4 13.24 0.4 ;
      RECT 3.01 -0.4 3.35 0.575 ;
      RECT 1.33 -0.4 3.01 0.4 ;
      RECT 0.99 -0.4 1.33 0.575 ;
      RECT 0 -0.4 0.99 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 21.385 4.64 22.44 5.44 ;
      RECT 21.045 4.085 21.385 5.44 ;
      RECT 20.125 4.64 21.045 5.44 ;
      RECT 19.785 4.085 20.125 5.44 ;
      RECT 18.79 4.64 19.785 5.44 ;
      RECT 18.385 4.465 18.79 5.44 ;
      RECT 14.09 4.64 18.385 5.44 ;
      RECT 13.75 4.01 14.09 5.44 ;
      RECT 12.65 4.64 13.75 5.44 ;
      RECT 12.31 4.01 12.65 5.44 ;
      RECT 3.66 4.64 12.31 5.44 ;
      RECT 3.32 3.765 3.66 5.44 ;
      RECT 1.445 4.64 3.32 5.44 ;
      RECT 1.105 4 1.445 5.44 ;
      RECT 0 4.64 1.105 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 21.02 2.21 21.25 3.835 ;
      RECT 17.265 3.605 21.02 3.835 ;
      RECT 20.075 1.005 20.305 2.43 ;
      RECT 19.055 1.005 20.075 1.235 ;
      RECT 18.59 1.495 19.45 1.725 ;
      RECT 18.59 3.125 19.365 3.355 ;
      RECT 18.825 0.63 19.055 1.235 ;
      RECT 15.91 0.63 18.825 0.86 ;
      RECT 18.36 1.09 18.59 3.355 ;
      RECT 16.49 1.09 18.36 1.32 ;
      RECT 18.165 2.305 18.36 2.67 ;
      RECT 17.93 1.55 18.13 1.78 ;
      RECT 17.93 3.03 17.985 3.37 ;
      RECT 17.7 1.55 17.93 3.37 ;
      RECT 17.645 3.03 17.7 3.37 ;
      RECT 17.21 1.55 17.405 1.78 ;
      RECT 17.21 3.295 17.265 4.105 ;
      RECT 16.98 1.55 17.21 4.105 ;
      RECT 16.925 3.295 16.98 4.105 ;
      RECT 16.49 3.155 16.545 3.965 ;
      RECT 16.26 1.09 16.49 3.965 ;
      RECT 16.205 3.155 16.26 3.965 ;
      RECT 15.68 0.63 15.91 3.35 ;
      RECT 15.66 3.12 15.68 3.35 ;
      RECT 15.375 3.12 15.66 4.095 ;
      RECT 15.165 0.635 15.395 2.88 ;
      RECT 15.32 3.275 15.375 4.095 ;
      RECT 15.15 0.635 15.165 1.035 ;
      RECT 12.745 0.805 15.15 1.035 ;
      RECT 14.755 1.405 14.935 3.05 ;
      RECT 14.755 3.44 14.81 4.26 ;
      RECT 14.705 1.405 14.755 4.26 ;
      RECT 14.34 1.405 14.705 1.635 ;
      RECT 14.525 2.82 14.705 4.26 ;
      RECT 14.47 3.44 14.525 4.26 ;
      RECT 14.245 1.92 14.475 2.29 ;
      RECT 13.37 3.46 14.47 3.69 ;
      RECT 14 1.35 14.34 1.69 ;
      RECT 13.26 1.92 14.245 2.15 ;
      RECT 13.03 3.46 13.37 4.305 ;
      RECT 13.03 1.265 13.26 2.15 ;
      RECT 12.195 1.265 13.03 1.495 ;
      RECT 12.195 3.46 13.03 3.69 ;
      RECT 12.195 1.725 12.78 1.955 ;
      RECT 12.515 0.66 12.745 1.035 ;
      RECT 9.705 0.66 12.515 0.89 ;
      RECT 11.965 1.13 12.195 1.495 ;
      RECT 11.965 1.725 12.195 3.78 ;
      RECT 10.165 1.13 11.965 1.36 ;
      RECT 11.505 1.595 11.735 4.295 ;
      RECT 10.395 1.595 11.505 1.825 ;
      RECT 9.97 4.065 11.505 4.295 ;
      RECT 11.035 2.06 11.265 3.82 ;
      RECT 10.165 2.06 11.035 2.29 ;
      RECT 7.185 3.59 11.035 3.82 ;
      RECT 10.58 3.1 10.785 3.33 ;
      RECT 10.35 2.525 10.58 3.33 ;
      RECT 9.705 2.525 10.35 2.755 ;
      RECT 9.935 1.13 10.165 2.29 ;
      RECT 9.685 4.065 9.97 4.41 ;
      RECT 9.475 0.63 9.705 2.755 ;
      RECT 4.395 4.18 9.685 4.41 ;
      RECT 9.19 3.095 9.48 3.325 ;
      RECT 8.285 0.63 9.475 0.86 ;
      RECT 8.96 1.26 9.19 3.325 ;
      RECT 8.72 1.26 8.96 1.49 ;
      RECT 7.65 3.095 8.96 3.325 ;
      RECT 8.285 2.635 8.72 2.865 ;
      RECT 8.055 0.63 8.285 2.865 ;
      RECT 7.565 1.23 7.65 3.325 ;
      RECT 7.42 0.63 7.565 3.325 ;
      RECT 7.335 0.63 7.42 1.46 ;
      RECT 6.12 0.63 7.335 0.86 ;
      RECT 6.955 1.875 7.185 3.86 ;
      RECT 6.845 1.875 6.955 2.105 ;
      RECT 5.045 3.63 6.955 3.86 ;
      RECT 6.615 1.13 6.845 2.105 ;
      RECT 6.41 3.04 6.52 3.38 ;
      RECT 6.18 2.4 6.41 3.38 ;
      RECT 6.12 2.4 6.18 2.63 ;
      RECT 5.89 0.63 6.12 2.63 ;
      RECT 3.815 0.63 5.89 0.86 ;
      RECT 5.59 3.045 5.82 3.385 ;
      RECT 5.48 1.09 5.59 3.385 ;
      RECT 5.36 1.09 5.48 3.33 ;
      RECT 4.28 1.09 5.36 1.32 ;
      RECT 5.275 1.55 5.36 1.92 ;
      RECT 4.815 2.505 5.045 3.86 ;
      RECT 4.775 2.505 4.815 2.735 ;
      RECT 4.545 1.55 4.775 2.735 ;
      RECT 4.165 3.295 4.395 4.41 ;
      RECT 4.05 1.09 4.28 1.555 ;
      RECT 4.025 3.295 4.165 3.58 ;
      RECT 3.78 1.325 4.05 1.555 ;
      RECT 3.78 3.295 4.025 3.525 ;
      RECT 3.585 0.63 3.815 1.04 ;
      RECT 3.55 1.325 3.78 3.525 ;
      RECT 0.52 0.81 3.585 1.04 ;
      RECT 2.79 1.325 3.55 1.555 ;
      RECT 2.95 3.295 3.55 3.525 ;
      RECT 2.93 2.09 3.27 2.43 ;
      RECT 2.58 3.295 2.95 3.58 ;
      RECT 2.035 2.145 2.93 2.375 ;
      RECT 2.45 1.27 2.79 1.61 ;
      RECT 1.965 4.055 2.4 4.285 ;
      RECT 2.035 1.46 2.09 1.8 ;
      RECT 1.84 1.46 2.035 2.375 ;
      RECT 1.735 3.45 1.965 4.285 ;
      RECT 1.805 1.46 1.84 3.08 ;
      RECT 1.75 1.46 1.805 1.8 ;
      RECT 1.61 2.145 1.805 3.08 ;
      RECT 0.52 3.45 1.735 3.68 ;
      RECT 1.5 2.74 1.61 3.08 ;
      RECT 0.465 0.81 0.52 1.55 ;
      RECT 0.465 2.83 0.52 4.25 ;
      RECT 0.29 0.81 0.465 4.25 ;
      RECT 0.235 1.21 0.29 4.25 ;
      RECT 0.18 1.21 0.235 1.55 ;
      RECT 0.18 2.83 0.235 4.25 ;
  END
END ADDFHX2

MACRO ADDFHX1
  CLASS CORE ;
  FOREIGN ADDFHX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.18 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ ADDFHXL ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.4991 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.544 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.945 1.845 14.965 2.075 ;
      RECT 14.715 1.37 14.945 3.52 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.6026 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.021 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.625 1.845 13.645 2.075 ;
      RECT 13.395 1.37 13.625 3.685 ;
      RECT 13.11 3.455 13.395 3.685 ;
     END
  END CO

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2988 ;
  ANTENNAPARTIALMETALAREA 0.2874 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5264 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.62 2.94 12.985 3.195 ;
      RECT 12.39 2.35 12.62 3.195 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.17 ;
  ANTENNAPARTIALMETALAREA 0.348 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.905 2.94 7.705 3.375 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4788 ;
  ANTENNAPARTIALMETALAREA 0.2515 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0971 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.715 1.845 1.105 2.49 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.44 -0.4 15.18 0.4 ;
      RECT 14.1 -0.4 14.44 0.575 ;
      RECT 13.085 -0.4 14.1 0.4 ;
      RECT 12.745 -0.4 13.085 0.575 ;
      RECT 7.655 -0.4 12.745 0.4 ;
      RECT 7.315 -0.4 7.655 0.575 ;
      RECT 1.76 -0.4 7.315 0.4 ;
      RECT 1.42 -0.4 1.76 0.575 ;
      RECT 0 -0.4 1.42 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.21 4.64 15.18 5.44 ;
      RECT 13.87 4.465 14.21 5.44 ;
      RECT 11.98 4.64 13.87 5.44 ;
      RECT 11.64 4.465 11.98 5.44 ;
      RECT 7.485 4.64 11.64 5.44 ;
      RECT 7.145 4.065 7.485 5.44 ;
      RECT 2.385 4.64 7.145 5.44 ;
      RECT 2.045 3.69 2.385 5.44 ;
      RECT 1.24 4.64 2.045 5.44 ;
      RECT 0.9 3.755 1.24 5.44 ;
      RECT 0 4.64 0.9 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 14.215 2.455 14.305 2.815 ;
      RECT 13.985 2.455 14.215 4.235 ;
      RECT 10.445 4.005 13.985 4.235 ;
      RECT 12.515 0.805 13.79 1.035 ;
      RECT 12.055 1.5 12.915 1.73 ;
      RECT 12.055 3.46 12.745 3.69 ;
      RECT 12.285 0.63 12.515 1.035 ;
      RECT 9.435 0.63 12.285 0.86 ;
      RECT 11.825 1.09 12.055 3.69 ;
      RECT 10.1 1.09 11.825 1.32 ;
      RECT 11.49 2.56 11.825 2.79 ;
      RECT 11.475 1.62 11.595 1.85 ;
      RECT 11.26 1.62 11.475 2.315 ;
      RECT 11.245 1.62 11.26 3.69 ;
      RECT 11.03 2.085 11.245 3.69 ;
      RECT 10.88 3.46 11.03 3.69 ;
      RECT 10.75 1.62 10.875 1.85 ;
      RECT 10.52 1.62 10.75 3.215 ;
      RECT 10.445 2.985 10.52 3.215 ;
      RECT 10.215 2.985 10.445 4.235 ;
      RECT 9.87 1.09 10.1 2.75 ;
      RECT 9.725 2.52 9.87 2.75 ;
      RECT 9.495 2.52 9.725 3.75 ;
      RECT 9.265 0.63 9.435 1.85 ;
      RECT 9.205 0.63 9.265 4.295 ;
      RECT 9.035 1.62 9.205 4.295 ;
      RECT 8.585 4.065 9.035 4.295 ;
      RECT 8.2 0.64 8.905 0.87 ;
      RECT 8.575 1.565 8.805 3.835 ;
      RECT 8.43 1.565 8.575 1.905 ;
      RECT 8.26 3.605 8.575 3.835 ;
      RECT 8.2 2.46 8.345 3.275 ;
      RECT 7.83 3.605 8.26 3.995 ;
      RECT 8.115 0.64 8.2 3.275 ;
      RECT 7.97 0.64 8.115 2.69 ;
      RECT 7.085 0.865 7.97 1.095 ;
      RECT 6.71 3.605 7.83 3.835 ;
      RECT 7.51 1.36 7.74 2.605 ;
      RECT 6.625 1.36 7.51 1.59 ;
      RECT 6.855 0.63 7.085 1.095 ;
      RECT 5.245 0.63 6.855 0.86 ;
      RECT 6.63 3.605 6.71 4.125 ;
      RECT 6.4 2.085 6.63 4.125 ;
      RECT 6.395 1.09 6.625 1.59 ;
      RECT 5.705 1.09 6.395 1.32 ;
      RECT 5.935 1.55 6.165 4.405 ;
      RECT 3.085 4.175 5.935 4.405 ;
      RECT 5.475 1.09 5.705 3.945 ;
      RECT 3.805 3.715 5.475 3.945 ;
      RECT 5.015 0.63 5.245 3.38 ;
      RECT 4.295 0.75 4.525 3.38 ;
      RECT 2.225 0.75 4.295 0.98 ;
      RECT 3.805 1.22 3.86 1.56 ;
      RECT 3.575 1.22 3.805 3.945 ;
      RECT 3.52 1.22 3.575 1.56 ;
      RECT 3.085 1.22 3.14 1.56 ;
      RECT 2.855 1.22 3.085 4.405 ;
      RECT 2.8 1.22 2.855 1.56 ;
      RECT 2.125 2.015 2.605 2.405 ;
      RECT 1.995 0.75 2.225 1.095 ;
      RECT 1.895 1.515 2.125 3.23 ;
      RECT 0.465 0.865 1.995 1.095 ;
      RECT 1.54 1.515 1.895 1.745 ;
      RECT 1.5 3 1.895 3.23 ;
      RECT 0.465 3.035 0.52 3.975 ;
      RECT 0.235 0.865 0.465 3.975 ;
      RECT 0.18 3.035 0.235 3.975 ;
  END
END ADDFHX1

#MACRO ANTENNA
#  CLASS CORE ;
#  FOREIGN ANTENNA 0 0 ;
#  ORIGIN 0 0 ;
#  SIZE 1.32 BY 5.04 ;
#  SYMMETRY X Y ;
#  SITE tsm3site ;
#
#  PIN A
#  DIRECTION INPUT ;
#  ANTENNADIFFAREA 1.0764 ;
#  ANTENNAPARTIALMETALAREA 0.3588 LAYER Metal1 ;
#  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
#     PORT
#      LAYER Metal1 ;
#      RECT 0.14 1.26 0.83 1.78 ;
#     END
#  END A
#
#  PIN VSS
#  DIRECTION INOUT ;
#  USE GROUND ;
#  SHAPE ABUTMENT ;
#     PORT
#      LAYER Metal1 ;
#      RECT 0 -0.4 1.32 0.4 ;
#     END
#  END VSS
#
#  PIN VDD
#  DIRECTION INOUT ;
#  USE POWER ;
#  SHAPE ABUTMENT ;
#     PORT
#      LAYER Metal1 ;
#      RECT 0 4.64 1.32 5.44 ;
#     END
#  END VDD
#END ANTENNA

MACRO RFRDX4
  CLASS CORE ;
  FOREIGN RFRDX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.96 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN RB
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0692 ;
  ANTENNADIFFAREA 0.4088 ;
  ANTENNAPARTIALMETALAREA 1.0377 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.823 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.665 1.46 3.775 1.845 ;
      RECT 3.44 1.46 3.665 2.075 ;
      RECT 3.435 1.46 3.44 2.1 ;
      RECT 3.3 1.845 3.435 2.1 ;
      RECT 3.3 2.635 3.35 3.08 ;
      RECT 3.07 1.845 3.3 3.08 ;
      RECT 1.64 1.845 3.07 2.075 ;
      RECT 3.01 2.635 3.07 3.08 ;
      RECT 1.41 1.845 1.64 2.53 ;
     END
  END RB

  PIN BRB
  DIRECTION OUTPUT ;
  ANTENNAGATEAREA 0.4704 ;
  ANTENNADIFFAREA 1.7454 ;
  ANTENNAPARTIALMETALAREA 1.5699 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.4802 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.41 3.135 2.75 3.475 ;
      RECT 1.535 3.19 2.41 3.42 ;
      RECT 1.355 2.855 1.535 3.42 ;
      RECT 1.18 2.855 1.355 3.76 ;
      RECT 1.18 0.78 1.285 1.615 ;
      RECT 1.175 0.78 1.18 1.845 ;
      RECT 1.175 2.38 1.18 3.78 ;
      RECT 0.945 0.78 1.175 3.78 ;
      RECT 0.8 2.38 0.945 3.78 ;
     END
  END BRB

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.045 -0.4 3.96 0.4 ;
      RECT 2.01 -0.4 2.045 0.575 ;
      RECT 1.67 -0.4 2.01 1.12 ;
      RECT 0.52 -0.4 1.67 0.4 ;
      RECT 0.52 0.78 0.56 1.12 ;
      RECT 0.22 -0.4 0.52 1.12 ;
      RECT 0.18 -0.4 0.22 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 2.16 4.64 3.96 5.44 ;
      RECT 1.82 3.94 2.16 5.44 ;
      RECT 0.56 4.64 1.82 5.44 ;
      RECT 0.22 3.94 0.56 5.44 ;
      RECT 0 4.64 0.22 5.44 ;
     END
  END VDD
END RFRDX4

MACRO RFRDX2
  CLASS CORE ;
  FOREIGN RFRDX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ RFRDX4 ;

  PIN RB
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5346 ;
  ANTENNADIFFAREA 0.4088 ;
  ANTENNAPARTIALMETALAREA 1.269 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.9201 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.03 0.97 3.08 1.31 ;
      RECT 2.8 0.97 3.03 3.655 ;
      RECT 2.74 0.97 2.8 1.31 ;
      RECT 1.105 1.845 2.8 2.075 ;
      RECT 2.69 3.195 2.8 3.655 ;
      RECT 0.875 1.845 1.105 2.6 ;
     END
  END RB

  PIN BRB
  DIRECTION OUTPUT ;
  ANTENNAGATEAREA 0.4788 ;
  ANTENNADIFFAREA 1.4964 ;
  ANTENNAPARTIALMETALAREA 1.1365 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.8866 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.065 2.785 2.405 3.125 ;
      RECT 1.765 2.84 2.065 3.125 ;
      RECT 0.56 2.84 1.765 3.07 ;
      RECT 0.445 1.46 0.56 1.845 ;
      RECT 0.52 2.84 0.56 3.655 ;
      RECT 0.445 2.635 0.52 3.655 ;
      RECT 0.215 1.46 0.445 3.655 ;
     END
  END BRB

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 -0.4 3.3 0.4 ;
      RECT 1.28 -0.4 1.32 0.575 ;
      RECT 0.94 -0.4 1.28 1.31 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.36 4.64 3.3 5.44 ;
      RECT 1.02 3.795 1.36 5.44 ;
      RECT 0 4.64 1.02 5.44 ;
     END
  END VDD
END RFRDX2

MACRO RFRDX1
  CLASS CORE ;
  FOREIGN RFRDX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.3 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ RFRDX4 ;

  PIN RB
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.27 ;
  ANTENNADIFFAREA 0.4088 ;
  ANTENNAPARTIALMETALAREA 1.383 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.3159 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.74 0.97 3.08 1.31 ;
      RECT 2.51 1.08 2.74 1.31 ;
      RECT 2.17 1.08 2.51 3.655 ;
      RECT 2.12 2.075 2.17 2.555 ;
      RECT 1.105 2.325 2.12 2.555 ;
      RECT 0.875 2.2 1.105 2.555 ;
     END
  END RB

  PIN BRB
  DIRECTION OUTPUT ;
  ANTENNAGATEAREA 0.4788 ;
  ANTENNADIFFAREA 0.756 ;
  ANTENNAPARTIALMETALAREA 1.0734 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.9449 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.855 2.785 1.91 3.125 ;
      RECT 1.57 2.785 1.855 3.195 ;
      RECT 0.56 2.965 1.57 3.195 ;
      RECT 0.33 0.97 0.56 3.655 ;
      RECT 0.22 0.97 0.33 1.31 ;
      RECT 0.22 3.195 0.33 3.655 ;
     END
  END BRB

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 -0.4 3.3 0.4 ;
      RECT 1.28 -0.4 1.32 0.575 ;
      RECT 0.94 -0.4 1.28 1.31 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 1.32 4.64 3.3 5.44 ;
      RECT 1.28 4.465 1.32 5.44 ;
      RECT 0.94 3.795 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
END RFRDX1

MACRO XOR3X4
  CLASS CORE ;
  FOREIGN XOR3X4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 19.8 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.467 ;
  ANTENNAPARTIALMETALAREA 1.1665 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.3089 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.95 2.94 19 4.34 ;
      RECT 18.9 0.955 18.95 4.34 ;
      RECT 18.72 0.835 18.9 4.34 ;
      RECT 18.56 0.835 18.72 1.645 ;
      RECT 18.62 2.74 18.72 4.34 ;
      RECT 18.6 2.74 18.62 3.08 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.1628 ;
  ANTENNAPARTIALMETALAREA 0.272 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4416 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.35 3.93 17.69 4.27 ;
      RECT 16.945 4.04 17.35 4.27 ;
      RECT 16.715 4.04 16.945 4.315 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.6604 ;
  ANTENNAPARTIALMETALAREA 0.5215 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2419 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12 2.675 12.11 3.015 ;
      RECT 11.77 1.575 12 3.015 ;
      RECT 11.52 1.575 11.77 2.1 ;
      RECT 11.435 1.845 11.52 2.1 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0884 ;
  ANTENNAPARTIALMETALAREA 0.2949 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.21 1.47 2.55 ;
      RECT 0.875 2.21 1.105 2.635 ;
      RECT 0.66 2.21 0.875 2.55 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.62 -0.4 19.8 0.4 ;
      RECT 19.28 -0.4 19.62 1.645 ;
      RECT 18.14 -0.4 19.28 0.4 ;
      RECT 17.8 -0.4 18.14 0.63 ;
      RECT 9.375 -0.4 17.8 0.4 ;
      RECT 9.035 -0.4 9.375 0.575 ;
      RECT 7.655 -0.4 9.035 0.4 ;
      RECT 7.315 -0.4 7.655 0.575 ;
      RECT 6.095 -0.4 7.315 0.4 ;
      RECT 5.755 -0.4 6.095 0.575 ;
      RECT 1.28 -0.4 5.755 0.4 ;
      RECT 0.94 -0.4 1.28 1.57 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.62 4.64 19.8 5.44 ;
      RECT 19.28 3.94 19.62 5.44 ;
      RECT 18.26 4.64 19.28 5.44 ;
      RECT 17.92 3.94 18.26 5.44 ;
      RECT 9.005 4.64 17.92 5.44 ;
      RECT 8.665 4.41 9.005 5.44 ;
      RECT 7.485 4.64 8.665 5.44 ;
      RECT 7.145 4.225 7.485 5.44 ;
      RECT 5.965 4.64 7.145 5.44 ;
      RECT 5.625 4.225 5.965 5.44 ;
      RECT 1.26 4.64 5.625 5.44 ;
      RECT 0.92 3.94 1.26 5.44 ;
      RECT 0 4.64 0.92 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 18.37 2.13 18.49 2.47 ;
      RECT 18.14 2.13 18.37 3.7 ;
      RECT 16.08 3.47 18.14 3.7 ;
      RECT 17.31 1.46 17.54 1.8 ;
      RECT 17.31 2.74 17.5 3.08 ;
      RECT 17.08 1.46 17.31 3.08 ;
      RECT 16.97 2.06 17.08 2.4 ;
      RECT 16.73 0.63 16.84 1.46 ;
      RECT 16.73 2.775 16.8 3.115 ;
      RECT 16.5 0.63 16.73 3.115 ;
      RECT 13.92 0.63 16.5 0.86 ;
      RECT 16.46 2.775 16.5 3.115 ;
      RECT 16.065 1.09 16.12 1.43 ;
      RECT 16.065 2.995 16.08 3.805 ;
      RECT 15.835 1.09 16.065 3.805 ;
      RECT 15.78 1.09 15.835 1.43 ;
      RECT 15.74 2.995 15.835 3.805 ;
      RECT 14.64 1.09 15.78 1.32 ;
      RECT 15.29 1.55 15.4 1.78 ;
      RECT 15.29 2.995 15.36 3.805 ;
      RECT 15.25 1.55 15.29 3.805 ;
      RECT 15.06 1.55 15.25 4.41 ;
      RECT 15.02 2.995 15.06 4.41 ;
      RECT 9.465 4.18 15.02 4.41 ;
      RECT 14.57 1.09 14.64 1.43 ;
      RECT 14.57 2.995 14.64 3.805 ;
      RECT 14.34 1.09 14.57 3.805 ;
      RECT 14.3 1.09 14.34 1.43 ;
      RECT 14.3 2.995 14.34 3.805 ;
      RECT 13.69 0.63 13.92 3.805 ;
      RECT 13.58 0.63 13.69 1.48 ;
      RECT 13.58 2.995 13.69 3.805 ;
      RECT 12.57 0.705 13.58 0.935 ;
      RECT 13.16 3.03 13.2 3.95 ;
      RECT 12.93 1.22 13.16 3.95 ;
      RECT 12.82 1.22 12.93 1.56 ;
      RECT 12.86 3.03 12.93 3.95 ;
      RECT 9.925 3.72 12.86 3.95 ;
      RECT 12.34 0.705 12.57 3.49 ;
      RECT 12.1 1.005 12.34 1.345 ;
      RECT 12.14 3.26 12.34 3.49 ;
      RECT 11.13 1.115 12.1 1.345 ;
      RECT 10.385 3.26 11.675 3.49 ;
      RECT 10.085 0.63 11.53 0.86 ;
      RECT 10.9 1.115 11.13 3.03 ;
      RECT 10.43 1.115 10.9 1.455 ;
      RECT 10.615 2.8 10.9 3.03 ;
      RECT 10.155 2.75 10.385 3.49 ;
      RECT 10.085 2.75 10.155 3.09 ;
      RECT 9.855 0.63 10.085 3.09 ;
      RECT 9.695 3.49 9.925 3.95 ;
      RECT 9.71 0.805 9.855 1.73 ;
      RECT 7.465 0.805 9.71 1.035 ;
      RECT 9.625 3.49 9.695 3.72 ;
      RECT 9.395 2 9.625 3.72 ;
      RECT 9.235 3.95 9.465 4.41 ;
      RECT 9.035 2 9.395 2.23 ;
      RECT 7.945 3.95 9.235 4.18 ;
      RECT 8.825 2.625 9.165 2.965 ;
      RECT 8.805 1.27 9.035 2.23 ;
      RECT 8.575 2.625 8.825 2.855 ;
      RECT 7.955 1.27 8.805 1.5 ;
      RECT 8.465 1.73 8.575 2.855 ;
      RECT 8.235 1.73 8.465 3.535 ;
      RECT 6.155 3.305 8.235 3.535 ;
      RECT 7.725 1.27 7.955 3.075 ;
      RECT 7.715 3.765 7.945 4.18 ;
      RECT 6.785 2.845 7.725 3.075 ;
      RECT 5.395 3.765 7.715 3.995 ;
      RECT 7.125 0.805 7.465 2.56 ;
      RECT 5.015 0.805 7.125 1.035 ;
      RECT 6.785 1.46 6.895 1.8 ;
      RECT 6.555 1.265 6.785 3.075 ;
      RECT 4.74 1.265 6.555 1.495 ;
      RECT 6.385 2.845 6.555 3.075 ;
      RECT 5.925 1.78 6.155 3.535 ;
      RECT 5.205 1.78 5.925 2.01 ;
      RECT 4.935 3.305 5.925 3.535 ;
      RECT 5.335 2.395 5.445 2.735 ;
      RECT 5.165 3.765 5.395 4.05 ;
      RECT 5.105 2.395 5.335 3.075 ;
      RECT 4.195 3.82 5.165 4.05 ;
      RECT 4.575 2.845 5.105 3.075 ;
      RECT 4.675 0.63 5.015 1.035 ;
      RECT 4.705 3.305 4.935 3.59 ;
      RECT 4.51 1.265 4.74 1.89 ;
      RECT 2.86 3.36 4.705 3.59 ;
      RECT 2.04 0.63 4.675 0.86 ;
      RECT 3.52 1.66 4.51 1.89 ;
      RECT 3.94 1.09 4.28 1.43 ;
      RECT 3.855 3.82 4.195 4.16 ;
      RECT 2.76 1.09 3.94 1.32 ;
      RECT 2.66 3.82 3.855 4.05 ;
      RECT 3.41 1.55 3.52 1.89 ;
      RECT 3.41 2.79 3.435 3.13 ;
      RECT 3.18 1.55 3.41 3.13 ;
      RECT 3.095 2.79 3.18 3.13 ;
      RECT 2.63 2.25 2.86 3.59 ;
      RECT 2.65 1.09 2.76 1.43 ;
      RECT 2.4 3.82 2.66 4.16 ;
      RECT 2.42 1.09 2.65 2.02 ;
      RECT 2.4 1.79 2.42 2.02 ;
      RECT 2.32 1.79 2.4 4.16 ;
      RECT 2.17 1.79 2.32 4.105 ;
      RECT 1.94 0.63 2.04 1.56 ;
      RECT 1.71 0.63 1.94 3.24 ;
      RECT 1.7 0.63 1.71 1.56 ;
      RECT 1.6 2.89 1.71 3.24 ;
      RECT 0.58 2.89 1.6 3.12 ;
      RECT 0.41 2.89 0.58 3.24 ;
      RECT 0.41 0.765 0.52 1.575 ;
      RECT 0.18 0.765 0.41 3.24 ;
  END
END XOR3X4

MACRO XOR3X2
  CLASS CORE ;
  FOREIGN XOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.88 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ XOR3X4 ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3572 ;
  ANTENNAPARTIALMETALAREA 0.718 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0846 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.7 0.955 11.75 3.025 ;
      RECT 11.665 0.835 11.7 3.08 ;
      RECT 11.52 0.835 11.665 3.195 ;
      RECT 11.36 0.835 11.52 1.645 ;
      RECT 11.435 2.74 11.52 3.195 ;
      RECT 11.36 2.74 11.435 3.08 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.2491 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.92 3.31 10.45 3.78 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 0.5353 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2472 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.025 2.405 7.045 2.635 ;
      RECT 6.915 2.405 7.025 3.23 ;
      RECT 6.685 1.79 6.915 3.23 ;
      RECT 6.365 1.79 6.685 2.13 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5442 ;
  ANTENNAPARTIALMETALAREA 0.2507 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.21 0.82 2.55 ;
      RECT 0.215 2.21 0.445 2.635 ;
      RECT 0.14 2.21 0.215 2.55 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.94 -0.4 11.88 0.4 ;
      RECT 10.6 -0.4 10.94 0.63 ;
      RECT 3.695 -0.4 10.6 0.4 ;
      RECT 3.355 -0.4 3.695 0.815 ;
      RECT 0.52 -0.4 3.355 0.4 ;
      RECT 0.18 -0.4 0.52 1.57 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.02 4.64 11.88 5.44 ;
      RECT 10.68 3.94 11.02 5.44 ;
      RECT 3.535 4.64 10.68 5.44 ;
      RECT 3.195 4.185 3.535 5.44 ;
      RECT 0.6 4.64 3.195 5.44 ;
      RECT 0.26 3.94 0.6 5.44 ;
      RECT 0 4.64 0.26 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 11.13 2.13 11.29 2.47 ;
      RECT 10.9 1 11.13 2.47 ;
      RECT 10.18 1 10.9 1.23 ;
      RECT 10.11 1.46 10.34 1.8 ;
      RECT 10.11 2.74 10.3 3.08 ;
      RECT 9.95 0.765 10.18 1.23 ;
      RECT 9.88 1.46 10.11 3.08 ;
      RECT 8.88 0.765 9.95 0.995 ;
      RECT 9.77 2.06 9.88 2.4 ;
      RECT 9.53 1.225 9.64 1.565 ;
      RECT 9.53 2.995 9.6 3.805 ;
      RECT 9.49 1.225 9.53 3.805 ;
      RECT 9.3 1.225 9.49 4.41 ;
      RECT 9.26 2.995 9.3 4.41 ;
      RECT 4.615 4.18 9.26 4.41 ;
      RECT 8.81 0.63 8.88 1.44 ;
      RECT 8.81 2.995 8.88 3.805 ;
      RECT 8.58 0.63 8.81 3.805 ;
      RECT 8.54 0.63 8.58 1.44 ;
      RECT 8.54 2.995 8.58 3.805 ;
      RECT 7.93 0.63 8.16 3.805 ;
      RECT 7.82 0.63 7.93 1.48 ;
      RECT 7.82 2.995 7.93 3.805 ;
      RECT 6.135 0.63 7.82 0.86 ;
      RECT 7.36 1.22 7.59 3.95 ;
      RECT 7.06 1.22 7.36 1.56 ;
      RECT 7.1 3.61 7.36 3.95 ;
      RECT 5.075 3.72 7.1 3.95 ;
      RECT 6.115 2.75 6.455 3.09 ;
      RECT 6.025 0.63 6.135 1.73 ;
      RECT 6.025 2.75 6.115 2.98 ;
      RECT 5.905 0.63 6.025 2.98 ;
      RECT 5.795 0.92 5.905 2.98 ;
      RECT 5.535 3.26 5.735 3.49 ;
      RECT 5.415 1.045 5.535 3.49 ;
      RECT 5.305 0.84 5.415 3.49 ;
      RECT 5.075 0.84 5.305 1.275 ;
      RECT 3.235 1.045 5.075 1.275 ;
      RECT 4.845 1.505 5.075 3.95 ;
      RECT 3.695 1.505 4.845 1.735 ;
      RECT 4.565 1.965 4.615 2.195 ;
      RECT 4.385 3.725 4.615 4.41 ;
      RECT 4.455 1.965 4.565 2.8 ;
      RECT 4.225 1.965 4.455 3.495 ;
      RECT 2 3.725 4.385 3.955 ;
      RECT 2.2 3.265 4.225 3.495 ;
      RECT 3.465 1.505 3.695 3.035 ;
      RECT 2.665 2.805 3.465 3.035 ;
      RECT 3.125 1.045 3.235 2.56 ;
      RECT 2.895 0.63 3.125 2.56 ;
      RECT 1.28 0.63 2.895 0.86 ;
      RECT 2.435 1.12 2.665 3.035 ;
      RECT 1.97 2.07 2.2 3.495 ;
      RECT 1.74 1.09 2 1.43 ;
      RECT 1.74 3.725 2 4.065 ;
      RECT 1.66 1.09 1.74 4.065 ;
      RECT 1.51 1.145 1.66 4.01 ;
      RECT 1.05 0.63 1.28 3.13 ;
      RECT 0.94 0.63 1.05 1.47 ;
      RECT 0.94 2.79 1.05 3.13 ;
  END
END XOR3X2

MACRO XNOR2X2_LVT
  CLASS CORE ;
  FOREIGN XNOR2X2_LVT 0 0 ;
  ORIGIN 0 0 ;
  SIZE 19.8 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.467 ;
  ANTENNAPARTIALMETALAREA 1.1665 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.3089 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.95 2.94 19 4.34 ;
      RECT 18.9 0.955 18.95 4.34 ;
      RECT 18.72 0.835 18.9 4.34 ;
      RECT 18.56 0.835 18.72 1.645 ;
      RECT 18.62 2.74 18.72 4.34 ;
      RECT 18.6 2.74 18.62 3.08 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.1628 ;
  ANTENNAPARTIALMETALAREA 0.272 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.4416 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.35 3.93 17.69 4.27 ;
      RECT 16.945 4.04 17.35 4.27 ;
      RECT 16.715 4.04 16.945 4.315 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.6604 ;
  ANTENNAPARTIALMETALAREA 0.5005 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.1995 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.96 2.675 12.07 3.015 ;
      RECT 11.73 1.575 11.96 3.015 ;
      RECT 11.52 1.575 11.73 2.1 ;
      RECT 11.435 1.845 11.52 2.1 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0884 ;
  ANTENNAPARTIALMETALAREA 0.2949 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.21 1.47 2.55 ;
      RECT 0.875 2.21 1.105 2.635 ;
      RECT 0.66 2.21 0.875 2.55 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.62 -0.4 19.8 0.4 ;
      RECT 19.28 -0.4 19.62 1.645 ;
      RECT 18.14 -0.4 19.28 0.4 ;
      RECT 17.8 -0.4 18.14 0.63 ;
      RECT 9.375 -0.4 17.8 0.4 ;
      RECT 9.035 -0.4 9.375 0.575 ;
      RECT 7.655 -0.4 9.035 0.4 ;
      RECT 7.315 -0.4 7.655 0.575 ;
      RECT 6.095 -0.4 7.315 0.4 ;
      RECT 5.755 -0.4 6.095 0.575 ;
      RECT 1.28 -0.4 5.755 0.4 ;
      RECT 0.94 -0.4 1.28 1.57 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 19.62 4.64 19.8 5.44 ;
      RECT 19.28 3.94 19.62 5.44 ;
      RECT 18.26 4.64 19.28 5.44 ;
      RECT 17.92 3.94 18.26 5.44 ;
      RECT 9.005 4.64 17.92 5.44 ;
      RECT 8.665 4.41 9.005 5.44 ;
      RECT 7.485 4.64 8.665 5.44 ;
      RECT 7.145 4.225 7.485 5.44 ;
      RECT 5.965 4.64 7.145 5.44 ;
      RECT 5.625 4.225 5.965 5.44 ;
      RECT 1.26 4.64 5.625 5.44 ;
      RECT 0.92 3.94 1.26 5.44 ;
      RECT 0 4.64 0.92 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 18.37 2.13 18.49 2.47 ;
      RECT 18.14 2.13 18.37 3.7 ;
      RECT 16.105 3.47 18.14 3.7 ;
      RECT 17.34 1.46 17.58 1.8 ;
      RECT 17.34 2.74 17.5 3.08 ;
      RECT 17.11 1.46 17.34 3.08 ;
      RECT 16.97 2.095 17.11 2.435 ;
      RECT 16.73 1.46 16.88 1.8 ;
      RECT 16.73 2.775 16.8 3.115 ;
      RECT 16.5 0.63 16.73 3.115 ;
      RECT 13.88 0.63 16.5 0.86 ;
      RECT 16.46 2.775 16.5 3.115 ;
      RECT 16.105 1.09 16.16 1.48 ;
      RECT 16.08 1.09 16.105 3.7 ;
      RECT 15.875 1.09 16.08 3.805 ;
      RECT 15.82 1.09 15.875 1.48 ;
      RECT 15.74 2.995 15.875 3.805 ;
      RECT 14.6 1.09 15.82 1.32 ;
      RECT 15.29 1.55 15.4 1.78 ;
      RECT 15.29 2.995 15.36 3.805 ;
      RECT 15.25 1.55 15.29 3.805 ;
      RECT 15.06 1.55 15.25 4.41 ;
      RECT 15.02 2.995 15.06 4.41 ;
      RECT 9.465 4.18 15.02 4.41 ;
      RECT 14.57 2.995 14.64 3.805 ;
      RECT 14.57 1.09 14.6 1.48 ;
      RECT 14.34 1.09 14.57 3.805 ;
      RECT 14.26 1.09 14.34 1.48 ;
      RECT 14.3 2.995 14.34 3.805 ;
      RECT 13.88 2.995 13.92 3.805 ;
      RECT 13.65 0.63 13.88 3.805 ;
      RECT 13.54 0.63 13.65 1.48 ;
      RECT 13.58 2.995 13.65 3.805 ;
      RECT 12.53 0.705 13.54 0.935 ;
      RECT 13.16 3.03 13.2 3.95 ;
      RECT 12.93 1.22 13.16 3.95 ;
      RECT 12.78 1.22 12.93 1.56 ;
      RECT 12.86 3.03 12.93 3.95 ;
      RECT 9.925 3.72 12.86 3.95 ;
      RECT 12.3 0.705 12.53 3.49 ;
      RECT 12.06 1.005 12.3 1.345 ;
      RECT 12.14 3.26 12.3 3.49 ;
      RECT 11.13 1.115 12.06 1.345 ;
      RECT 10.385 3.26 11.675 3.49 ;
      RECT 10.085 0.63 11.49 0.86 ;
      RECT 10.9 1.115 11.13 3.03 ;
      RECT 10.39 1.115 10.9 1.455 ;
      RECT 10.615 2.8 10.9 3.03 ;
      RECT 10.155 2.745 10.385 3.49 ;
      RECT 10.085 2.745 10.155 3.085 ;
      RECT 9.855 0.63 10.085 3.085 ;
      RECT 9.695 3.49 9.925 3.95 ;
      RECT 9.67 0.805 9.855 1.73 ;
      RECT 9.625 3.49 9.695 3.72 ;
      RECT 7.465 0.805 9.67 1.035 ;
      RECT 9.395 2 9.625 3.72 ;
      RECT 9.235 3.95 9.465 4.41 ;
      RECT 9.035 2 9.395 2.23 ;
      RECT 7.945 3.95 9.235 4.18 ;
      RECT 8.825 2.625 9.165 2.965 ;
      RECT 8.805 1.27 9.035 2.23 ;
      RECT 8.575 2.625 8.825 2.855 ;
      RECT 7.955 1.27 8.805 1.5 ;
      RECT 8.465 1.73 8.575 2.855 ;
      RECT 8.235 1.73 8.465 3.535 ;
      RECT 6.155 3.305 8.235 3.535 ;
      RECT 7.725 1.27 7.955 3.075 ;
      RECT 7.715 3.765 7.945 4.18 ;
      RECT 6.785 2.845 7.725 3.075 ;
      RECT 5.395 3.765 7.715 3.995 ;
      RECT 7.125 0.805 7.465 2.56 ;
      RECT 5.015 0.805 7.125 1.035 ;
      RECT 6.785 1.46 6.895 1.8 ;
      RECT 6.555 1.265 6.785 3.075 ;
      RECT 4.74 1.265 6.555 1.495 ;
      RECT 6.385 2.845 6.555 3.075 ;
      RECT 5.925 1.725 6.155 3.535 ;
      RECT 5.205 1.725 5.925 2.065 ;
      RECT 4.935 3.305 5.925 3.535 ;
      RECT 5.335 2.395 5.445 2.735 ;
      RECT 5.165 3.765 5.395 4.105 ;
      RECT 5.105 2.395 5.335 3.075 ;
      RECT 4.195 3.875 5.165 4.105 ;
      RECT 4.575 2.845 5.105 3.075 ;
      RECT 4.675 0.63 5.015 1.035 ;
      RECT 4.705 3.305 4.935 3.59 ;
      RECT 4.51 1.265 4.74 1.89 ;
      RECT 2.86 3.36 4.705 3.59 ;
      RECT 2.04 0.63 4.675 0.86 ;
      RECT 3.52 1.66 4.51 1.89 ;
      RECT 3.94 1.09 4.28 1.43 ;
      RECT 3.855 3.82 4.195 4.16 ;
      RECT 2.76 1.09 3.94 1.32 ;
      RECT 2.66 3.82 3.855 4.05 ;
      RECT 3.41 1.55 3.52 1.89 ;
      RECT 3.41 2.79 3.435 3.13 ;
      RECT 3.18 1.55 3.41 3.13 ;
      RECT 3.095 2.79 3.18 3.13 ;
      RECT 2.63 2.25 2.86 3.59 ;
      RECT 2.65 1.09 2.76 1.43 ;
      RECT 2.4 3.82 2.66 4.16 ;
      RECT 2.42 1.09 2.65 2.02 ;
      RECT 2.4 1.79 2.42 2.02 ;
      RECT 2.32 1.79 2.4 4.16 ;
      RECT 2.17 1.79 2.32 4.105 ;
      RECT 1.94 0.63 2.04 1.56 ;
      RECT 1.71 0.63 1.94 3.24 ;
      RECT 1.7 0.63 1.71 1.56 ;
      RECT 1.6 2.89 1.71 3.24 ;
      RECT 0.58 2.89 1.6 3.12 ;
      RECT 0.41 2.89 0.58 3.24 ;
      RECT 0.41 0.765 0.52 1.575 ;
      RECT 0.18 0.765 0.41 3.24 ;
  END
END XNOR2X2_LVT

MACRO XNOR3X2
  CLASS CORE ;
  FOREIGN XNOR3X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.88 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ XNOR2X2_LVT ;

  PIN Y
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3572 ;
  ANTENNAPARTIALMETALAREA 0.718 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0846 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.7 0.955 11.75 3.025 ;
      RECT 11.665 0.835 11.7 3.08 ;
      RECT 11.52 0.835 11.665 3.195 ;
      RECT 11.36 0.835 11.52 1.645 ;
      RECT 11.435 2.74 11.52 3.195 ;
      RECT 11.36 2.74 11.435 3.08 ;
     END
  END Y

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.2491 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.06 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.92 3.31 10.45 3.78 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 0.5353 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2472 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.025 2.405 7.045 2.635 ;
      RECT 6.915 2.405 7.025 3.23 ;
      RECT 6.685 1.79 6.915 3.23 ;
      RECT 6.365 1.79 6.685 2.13 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5442 ;
  ANTENNAPARTIALMETALAREA 0.2507 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1713 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.21 0.82 2.55 ;
      RECT 0.215 2.21 0.445 2.635 ;
      RECT 0.14 2.21 0.215 2.55 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 10.94 -0.4 11.88 0.4 ;
      RECT 10.6 -0.4 10.94 0.63 ;
      RECT 3.695 -0.4 10.6 0.4 ;
      RECT 3.355 -0.4 3.695 0.815 ;
      RECT 0.52 -0.4 3.355 0.4 ;
      RECT 0.18 -0.4 0.52 1.57 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.02 4.64 11.88 5.44 ;
      RECT 10.68 3.94 11.02 5.44 ;
      RECT 3.535 4.64 10.68 5.44 ;
      RECT 3.195 4.185 3.535 5.44 ;
      RECT 0.6 4.64 3.195 5.44 ;
      RECT 0.26 3.94 0.6 5.44 ;
      RECT 0 4.64 0.26 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 11.13 2.13 11.29 2.47 ;
      RECT 10.9 1 11.13 2.47 ;
      RECT 10.18 1 10.9 1.23 ;
      RECT 10.11 1.46 10.34 1.8 ;
      RECT 10.11 2.74 10.3 3.08 ;
      RECT 9.95 0.63 10.18 1.23 ;
      RECT 9.88 1.46 10.11 3.08 ;
      RECT 8.88 0.63 9.95 0.86 ;
      RECT 9.77 2.21 9.88 2.55 ;
      RECT 9.53 1.14 9.64 1.48 ;
      RECT 9.53 2.995 9.6 3.805 ;
      RECT 9.49 1.14 9.53 3.805 ;
      RECT 9.3 1.14 9.49 4.41 ;
      RECT 9.26 2.995 9.3 4.41 ;
      RECT 4.615 4.18 9.26 4.41 ;
      RECT 8.81 0.63 8.88 1.44 ;
      RECT 8.81 2.995 8.88 3.805 ;
      RECT 8.58 0.63 8.81 3.805 ;
      RECT 8.54 0.63 8.58 1.44 ;
      RECT 8.54 2.995 8.58 3.805 ;
      RECT 7.93 0.63 8.16 3.805 ;
      RECT 7.82 0.63 7.93 1.48 ;
      RECT 7.82 2.995 7.93 3.805 ;
      RECT 6.135 0.63 7.82 0.86 ;
      RECT 7.36 1.22 7.59 3.95 ;
      RECT 7.06 1.22 7.36 1.56 ;
      RECT 7.1 3.61 7.36 3.95 ;
      RECT 5.075 3.72 7.1 3.95 ;
      RECT 6.115 2.75 6.455 3.09 ;
      RECT 6.025 0.63 6.135 1.73 ;
      RECT 6.025 2.75 6.115 2.98 ;
      RECT 5.905 0.63 6.025 2.98 ;
      RECT 5.795 0.92 5.905 2.98 ;
      RECT 5.535 3.26 5.735 3.49 ;
      RECT 5.415 1.045 5.535 3.49 ;
      RECT 5.305 0.84 5.415 3.49 ;
      RECT 5.075 0.84 5.305 1.275 ;
      RECT 3.235 1.045 5.075 1.275 ;
      RECT 4.845 1.505 5.075 3.95 ;
      RECT 3.695 1.505 4.845 1.735 ;
      RECT 4.565 1.965 4.615 2.195 ;
      RECT 4.385 3.725 4.615 4.41 ;
      RECT 4.455 1.965 4.565 2.8 ;
      RECT 4.225 1.965 4.455 3.495 ;
      RECT 2 3.725 4.385 3.955 ;
      RECT 2.2 3.265 4.225 3.495 ;
      RECT 3.465 1.505 3.695 3.035 ;
      RECT 2.665 2.805 3.465 3.035 ;
      RECT 3.125 1.045 3.235 2.56 ;
      RECT 2.895 0.63 3.125 2.56 ;
      RECT 1.28 0.63 2.895 0.86 ;
      RECT 2.435 1.12 2.665 3.035 ;
      RECT 1.97 2.07 2.2 3.495 ;
      RECT 1.74 1.09 2 1.43 ;
      RECT 1.74 3.725 2 4.065 ;
      RECT 1.66 1.09 1.74 4.065 ;
      RECT 1.51 1.145 1.66 4.01 ;
      RECT 1.05 0.63 1.28 3.13 ;
      RECT 0.94 0.63 1.05 1.47 ;
      RECT 0.94 2.79 1.05 3.13 ;
  END
END XNOR3X2

MACRO AFCSHCONX4
  CLASS CORE ;
  FOREIGN AFCSHCONX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 31.02 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 1.1475 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1552 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 30.88 0.97 30.89 3.025 ;
      RECT 30.66 0.97 30.88 4.34 ;
      RECT 30.5 0.97 30.66 1.78 ;
      RECT 30.5 2.74 30.66 4.34 ;
     END
  END S

  PIN CS
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.44 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0935 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 29.81 1.26 30.22 1.54 ;
      RECT 29.58 1.26 29.81 2.43 ;
      RECT 29.415 2.09 29.58 2.43 ;
     END
  END CS

  PIN CO1N
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.522 ;
  ANTENNAPARTIALMETALAREA 2.1685 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.3386 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.02 2.205 20.38 2.435 ;
      RECT 17.02 3.685 20.38 3.915 ;
      RECT 16.735 2.205 17.02 3.915 ;
      RECT 16.715 2.38 16.735 3.915 ;
      RECT 16.64 2.38 16.715 3.78 ;
     END
  END CO1N

  PIN CO0N
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.513 ;
  ANTENNAPARTIALMETALAREA 2.1583 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.2326 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.315 2.38 16.36 3.78 ;
      RECT 15.98 2.205 16.315 3.915 ;
      RECT 12.67 2.205 15.98 2.435 ;
      RECT 12.67 3.685 15.98 3.915 ;
     END
  END CO0N

  PIN CI1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0194 ;
  ANTENNAPARTIALMETALAREA 0.2227 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0017 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 24.56 2.28 25.055 2.73 ;
     END
  END CI1

  PIN CI0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0068 ;
  ANTENNAPARTIALMETALAREA 0.2296 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.88 2.25 8.44 2.66 ;
     END
  END CI0

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.4493 ;
  ANTENNAPARTIALMETALAREA 0.252 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1289 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.41 4.03 7.12 4.385 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.759 ;
  ANTENNAPARTIALMETALAREA 0.2881 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5158 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.105 1.18 2.445 ;
      RECT 0.875 2.105 1.105 3.195 ;
      RECT 0.84 2.105 0.875 2.445 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 30.08 -0.4 31.02 0.4 ;
      RECT 29.74 -0.4 30.08 0.63 ;
      RECT 28.55 -0.4 29.74 0.4 ;
      RECT 28.21 -0.4 28.55 1.78 ;
      RECT 25.375 -0.4 28.21 0.4 ;
      RECT 25.035 -0.4 25.375 0.575 ;
      RECT 24.015 -0.4 25.035 0.4 ;
      RECT 23.675 -0.4 24.015 0.575 ;
      RECT 9.375 -0.4 23.675 0.4 ;
      RECT 9.035 -0.4 9.375 0.575 ;
      RECT 8.015 -0.4 9.035 0.4 ;
      RECT 7.675 -0.4 8.015 0.575 ;
      RECT 2.38 -0.4 7.675 0.4 ;
      RECT 2.04 -0.4 2.38 0.63 ;
      RECT 1.2 -0.4 2.04 0.4 ;
      RECT 0.86 -0.4 1.2 0.63 ;
      RECT 0 -0.4 0.86 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 30.16 4.64 31.02 5.44 ;
      RECT 29.82 3.94 30.16 5.44 ;
      RECT 29.215 4.64 29.82 5.44 ;
      RECT 28.875 3.76 29.215 5.44 ;
      RECT 25.375 4.64 28.875 5.44 ;
      RECT 25.035 4.465 25.375 5.44 ;
      RECT 24.015 4.64 25.035 5.44 ;
      RECT 23.675 4.465 24.015 5.44 ;
      RECT 9.375 4.64 23.675 5.44 ;
      RECT 9.035 4.465 9.375 5.44 ;
      RECT 8.015 4.64 9.035 5.44 ;
      RECT 7.675 4.465 8.015 5.44 ;
      RECT 2.42 4.64 7.675 5.44 ;
      RECT 2.08 3.94 2.42 5.44 ;
      RECT 1.16 4.64 2.08 5.44 ;
      RECT 0.82 4.09 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 30.27 2.17 30.43 2.51 ;
      RECT 30.04 2.17 30.27 3.505 ;
      RECT 28.64 3.275 30.04 3.505 ;
      RECT 29.18 1.46 29.345 1.8 ;
      RECT 29.18 2.795 29.345 3.025 ;
      RECT 28.95 1.46 29.18 3.025 ;
      RECT 28.18 2.795 28.95 3.025 ;
      RECT 28.41 3.275 28.64 4.405 ;
      RECT 26.8 4.175 28.41 4.405 ;
      RECT 27.95 2.795 28.18 3.93 ;
      RECT 27.98 2.095 28.09 2.325 ;
      RECT 27.75 0.815 27.98 2.325 ;
      RECT 27.26 3.7 27.95 3.93 ;
      RECT 22.12 0.815 27.75 1.045 ;
      RECT 27.52 2.62 27.72 3.45 ;
      RECT 27.49 1.38 27.52 3.45 ;
      RECT 27.29 1.38 27.49 2.85 ;
      RECT 27.06 3.08 27.26 3.93 ;
      RECT 27.03 2.17 27.06 3.93 ;
      RECT 26.83 2.17 27.03 3.31 ;
      RECT 26.595 1.38 26.855 1.72 ;
      RECT 26.595 3.54 26.8 4.405 ;
      RECT 26.57 1.38 26.595 4.405 ;
      RECT 26.365 1.38 26.57 3.77 ;
      RECT 25.905 1.38 26.135 3.965 ;
      RECT 25.795 1.38 25.905 1.72 ;
      RECT 25.795 3.155 25.905 3.965 ;
      RECT 25.515 2.39 25.625 2.73 ;
      RECT 25.285 1.275 25.515 2.73 ;
      RECT 22.64 1.275 25.285 1.505 ;
      RECT 24.325 1.735 24.695 1.965 ;
      RECT 24.32 2.96 24.64 3.775 ;
      RECT 24.32 1.735 24.325 2.665 ;
      RECT 24.09 1.735 24.32 3.775 ;
      RECT 23.395 2.435 24.09 2.665 ;
      RECT 21.635 3.545 24.09 3.775 ;
      RECT 23.125 3.08 23.305 3.31 ;
      RECT 23.125 1.735 23.255 1.965 ;
      RECT 22.895 1.735 23.125 3.31 ;
      RECT 22.41 1.275 22.64 3.31 ;
      RECT 22.195 1.735 22.41 1.965 ;
      RECT 22.245 3.08 22.41 3.31 ;
      RECT 21.89 0.815 22.12 1.485 ;
      RECT 20.965 1.255 21.89 1.485 ;
      RECT 21.635 1.735 21.76 1.965 ;
      RECT 21.405 1.735 21.635 3.775 ;
      RECT 10.09 0.735 21.465 0.965 ;
      RECT 17.43 2.965 21.405 3.195 ;
      RECT 12.285 4.18 21.295 4.41 ;
      RECT 20.735 1.255 20.965 1.965 ;
      RECT 10.84 1.735 20.735 1.965 ;
      RECT 7.28 1.275 20.38 1.505 ;
      RECT 11.975 2.965 15.62 3.195 ;
      RECT 11.755 4.005 12.285 4.41 ;
      RECT 11.975 2.195 12.085 2.425 ;
      RECT 11.745 2.195 11.975 3.775 ;
      RECT 7.95 4.005 11.755 4.235 ;
      RECT 8.915 3.545 11.745 3.775 ;
      RECT 10.61 1.735 10.84 3.31 ;
      RECT 10.515 1.735 10.61 1.965 ;
      RECT 10.465 3.08 10.61 3.31 ;
      RECT 9.925 1.735 10.155 3.31 ;
      RECT 9.86 0.735 10.09 1.045 ;
      RECT 9.795 1.735 9.925 1.965 ;
      RECT 9.745 3.08 9.925 3.31 ;
      RECT 7.28 0.815 9.86 1.045 ;
      RECT 8.915 2.435 9.655 2.665 ;
      RECT 8.685 1.735 8.915 3.775 ;
      RECT 8.355 1.735 8.685 1.965 ;
      RECT 8.41 2.95 8.685 3.775 ;
      RECT 7.72 3.57 7.95 4.235 ;
      RECT 6.625 3.57 7.72 3.8 ;
      RECT 7.28 3.045 7.335 3.275 ;
      RECT 7.05 0.63 7.28 1.045 ;
      RECT 7.05 1.275 7.28 3.275 ;
      RECT 5.245 0.63 7.05 0.86 ;
      RECT 6.855 2.47 7.05 3.275 ;
      RECT 6.625 1.09 6.745 2.24 ;
      RECT 6.515 1.09 6.625 3.8 ;
      RECT 5.705 1.09 6.515 1.32 ;
      RECT 6.395 2.01 6.515 3.8 ;
      RECT 6.165 1.55 6.275 1.78 ;
      RECT 5.935 1.55 6.165 4.405 ;
      RECT 3.1 4.175 5.935 4.405 ;
      RECT 5.475 1.09 5.705 3.945 ;
      RECT 3.86 3.715 5.475 3.945 ;
      RECT 5.015 0.63 5.245 3.485 ;
      RECT 4.47 1.075 4.58 1.415 ;
      RECT 4.47 3.145 4.58 3.485 ;
      RECT 4.24 0.63 4.47 3.485 ;
      RECT 3.1 0.63 4.24 0.86 ;
      RECT 3.805 1.22 3.86 1.56 ;
      RECT 3.805 3.135 3.86 3.945 ;
      RECT 3.575 1.22 3.805 3.945 ;
      RECT 3.52 1.22 3.575 1.56 ;
      RECT 3.52 3.135 3.575 3.945 ;
      RECT 3.1 1.325 3.14 1.665 ;
      RECT 2.87 0.63 3.1 1.095 ;
      RECT 2.87 1.325 3.1 4.405 ;
      RECT 0.52 0.865 2.87 1.095 ;
      RECT 2.8 1.325 2.87 1.665 ;
      RECT 2.76 2.74 2.87 3.08 ;
      RECT 1.84 2.04 2.585 2.38 ;
      RECT 1.61 1.46 1.84 3.08 ;
      RECT 1.5 1.46 1.61 1.8 ;
      RECT 1.5 2.74 1.61 3.08 ;
      RECT 0.29 0.865 0.52 3.08 ;
      RECT 0.18 1.46 0.29 1.8 ;
      RECT 0.18 2.74 0.29 3.08 ;
  END
END AFCSHCONX4

MACRO AFCSHCONX2
  CLASS CORE ;
  FOREIGN AFCSHCONX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 28.38 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AFCSHCONX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 1.1475 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1552 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 28.24 0.97 28.25 3.025 ;
      RECT 28.02 0.97 28.24 4.34 ;
      RECT 27.86 0.97 28.02 1.78 ;
      RECT 27.86 2.74 28.02 4.34 ;
     END
  END S

  PIN CS
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.44 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0935 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 27.17 1.26 27.58 1.54 ;
      RECT 26.94 1.26 27.17 2.43 ;
      RECT 26.775 2.09 26.94 2.43 ;
     END
  END CS

  PIN CO1N
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.3194 ;
  ANTENNAPARTIALMETALAREA 1.1931 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.3212 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.68 3.48 18.415 3.71 ;
      RECT 17.68 2.2 18.195 2.43 ;
      RECT 17.45 2.2 17.68 3.78 ;
      RECT 17.3 2.94 17.45 3.78 ;
      RECT 16.3 3.48 17.3 3.71 ;
      RECT 16.07 3.135 16.3 3.945 ;
     END
  END CO1N

  PIN CO0N
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.3194 ;
  ANTENNAPARTIALMETALAREA 1.1552 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.1463 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.23 3.135 14.46 3.945 ;
      RECT 13.06 3.48 14.23 3.71 ;
      RECT 12.91 2.94 13.06 3.78 ;
      RECT 12.68 2.195 12.91 3.78 ;
      RECT 12.335 2.195 12.68 2.425 ;
      RECT 12.115 3.48 12.68 3.71 ;
     END
  END CO0N

  PIN CI1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4791 ;
  ANTENNAPARTIALMETALAREA 0.2295 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.415 2.39 22.435 2.73 ;
      RECT 21.92 2.28 22.415 2.73 ;
     END
  END CI1

  PIN CI0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4818 ;
  ANTENNAPARTIALMETALAREA 0.2296 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.88 2.25 8.44 2.66 ;
     END
  END CI0

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.4493 ;
  ANTENNAPARTIALMETALAREA 0.252 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1289 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.41 4.03 7.12 4.385 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.759 ;
  ANTENNAPARTIALMETALAREA 0.2881 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5158 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.105 1.18 2.445 ;
      RECT 0.875 2.105 1.105 3.195 ;
      RECT 0.84 2.105 0.875 2.445 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 27.44 -0.4 28.38 0.4 ;
      RECT 27.1 -0.4 27.44 0.63 ;
      RECT 25.92 -0.4 27.1 0.4 ;
      RECT 25.69 -0.4 25.92 1.78 ;
      RECT 22.855 -0.4 25.69 0.4 ;
      RECT 22.515 -0.4 22.855 0.575 ;
      RECT 21.425 -0.4 22.515 0.4 ;
      RECT 21.085 -0.4 21.425 0.575 ;
      RECT 9.445 -0.4 21.085 0.4 ;
      RECT 9.105 -0.4 9.445 0.575 ;
      RECT 8.015 -0.4 9.105 0.4 ;
      RECT 7.675 -0.4 8.015 0.575 ;
      RECT 2.38 -0.4 7.675 0.4 ;
      RECT 2.04 -0.4 2.38 0.63 ;
      RECT 1.2 -0.4 2.04 0.4 ;
      RECT 0.86 -0.4 1.2 0.63 ;
      RECT 0 -0.4 0.86 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 27.52 4.64 28.38 5.44 ;
      RECT 27.18 3.94 27.52 5.44 ;
      RECT 26.695 4.64 27.18 5.44 ;
      RECT 26.355 3.76 26.695 5.44 ;
      RECT 22.855 4.64 26.355 5.44 ;
      RECT 22.515 4.465 22.855 5.44 ;
      RECT 21.475 4.64 22.515 5.44 ;
      RECT 21.135 4.465 21.475 5.44 ;
      RECT 9.395 4.64 21.135 5.44 ;
      RECT 9.055 4.465 9.395 5.44 ;
      RECT 8.015 4.64 9.055 5.44 ;
      RECT 7.675 4.465 8.015 5.44 ;
      RECT 2.42 4.64 7.675 5.44 ;
      RECT 2.08 3.94 2.42 5.44 ;
      RECT 1.16 4.64 2.08 5.44 ;
      RECT 0.82 4.09 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 27.63 2.17 27.79 2.51 ;
      RECT 27.4 2.17 27.63 3.505 ;
      RECT 26.12 3.275 27.4 3.505 ;
      RECT 26.53 1.46 26.695 1.8 ;
      RECT 26.53 2.795 26.695 3.025 ;
      RECT 26.3 1.46 26.53 3.025 ;
      RECT 25.66 2.795 26.3 3.025 ;
      RECT 25.89 3.275 26.12 4.405 ;
      RECT 24.28 4.175 25.89 4.405 ;
      RECT 25.43 2.795 25.66 3.915 ;
      RECT 25.46 2.095 25.57 2.325 ;
      RECT 25.23 0.815 25.46 2.325 ;
      RECT 24.74 3.685 25.43 3.915 ;
      RECT 19.67 0.815 25.23 1.045 ;
      RECT 25 2.62 25.2 3.45 ;
      RECT 24.97 1.38 25 3.45 ;
      RECT 24.77 1.38 24.97 2.85 ;
      RECT 24.54 3.08 24.74 3.915 ;
      RECT 24.51 2.17 24.54 3.915 ;
      RECT 24.31 2.17 24.51 3.31 ;
      RECT 24.075 1.38 24.335 1.72 ;
      RECT 24.075 3.54 24.28 4.405 ;
      RECT 24.05 1.38 24.075 4.405 ;
      RECT 23.845 1.38 24.05 3.77 ;
      RECT 23.385 1.38 23.615 3.965 ;
      RECT 23.275 1.38 23.385 1.72 ;
      RECT 23.275 3.155 23.385 3.965 ;
      RECT 22.995 2.39 23.105 2.73 ;
      RECT 22.765 1.275 22.995 2.73 ;
      RECT 20.195 1.275 22.765 1.505 ;
      RECT 21.69 1.735 22.175 1.965 ;
      RECT 21.69 2.96 22.12 3.8 ;
      RECT 21.46 1.735 21.69 3.8 ;
      RECT 21.005 2.435 21.46 2.665 ;
      RECT 19.38 3.57 21.46 3.8 ;
      RECT 20.735 3.08 20.915 3.31 ;
      RECT 20.735 1.735 20.865 1.965 ;
      RECT 20.505 1.735 20.735 3.31 ;
      RECT 19.965 1.275 20.195 3.31 ;
      RECT 19.335 1.735 19.965 1.965 ;
      RECT 19.855 3.08 19.965 3.31 ;
      RECT 19.44 0.815 19.67 1.485 ;
      RECT 18.135 1.255 19.44 1.485 ;
      RECT 19.15 2.2 19.38 4.4 ;
      RECT 18.575 2.2 19.15 2.43 ;
      RECT 10.09 0.735 18.96 0.965 ;
      RECT 17.905 1.255 18.135 1.965 ;
      RECT 15.84 1.735 17.905 1.965 ;
      RECT 15.38 1.275 17.435 1.505 ;
      RECT 10.075 4.18 16.71 4.41 ;
      RECT 15.61 1.735 15.84 3.5 ;
      RECT 14.92 3.27 15.61 3.5 ;
      RECT 15.15 1.275 15.38 3.035 ;
      RECT 7.28 1.275 15.15 1.505 ;
      RECT 14.69 1.735 14.92 3.5 ;
      RECT 10.71 1.735 14.69 1.965 ;
      RECT 11.47 2.195 11.955 2.425 ;
      RECT 11.24 2.195 11.47 3.945 ;
      RECT 11.095 3.545 11.24 3.945 ;
      RECT 8.915 3.545 11.095 3.775 ;
      RECT 10.48 1.735 10.71 3.31 ;
      RECT 10.385 1.735 10.48 1.965 ;
      RECT 10.335 3.08 10.48 3.31 ;
      RECT 9.86 0.735 10.09 1.045 ;
      RECT 9.845 4.005 10.075 4.41 ;
      RECT 9.795 1.735 10.025 3.31 ;
      RECT 7.28 0.815 9.86 1.045 ;
      RECT 7.95 4.005 9.845 4.235 ;
      RECT 9.665 1.735 9.795 1.965 ;
      RECT 9.615 3.08 9.795 3.31 ;
      RECT 8.915 2.435 9.525 2.665 ;
      RECT 8.685 1.735 8.915 3.775 ;
      RECT 8.355 1.735 8.685 1.965 ;
      RECT 8.41 2.95 8.685 3.775 ;
      RECT 7.72 3.57 7.95 4.235 ;
      RECT 6.625 3.57 7.72 3.8 ;
      RECT 7.28 3.045 7.335 3.275 ;
      RECT 7.05 0.63 7.28 1.045 ;
      RECT 7.05 1.275 7.28 3.275 ;
      RECT 5.245 0.63 7.05 0.86 ;
      RECT 6.855 2.47 7.05 3.275 ;
      RECT 6.625 1.09 6.745 2.24 ;
      RECT 6.515 1.09 6.625 3.8 ;
      RECT 5.705 1.09 6.515 1.32 ;
      RECT 6.395 2.01 6.515 3.8 ;
      RECT 6.165 1.55 6.275 1.78 ;
      RECT 5.935 1.55 6.165 4.405 ;
      RECT 3.1 4.175 5.935 4.405 ;
      RECT 5.475 1.09 5.705 3.945 ;
      RECT 3.86 3.715 5.475 3.945 ;
      RECT 5.015 0.63 5.245 3.485 ;
      RECT 4.47 1.075 4.58 1.415 ;
      RECT 4.47 3.145 4.58 3.485 ;
      RECT 4.24 0.63 4.47 3.485 ;
      RECT 3.1 0.63 4.24 0.86 ;
      RECT 3.805 1.22 3.86 1.56 ;
      RECT 3.805 3.135 3.86 3.945 ;
      RECT 3.575 1.22 3.805 3.945 ;
      RECT 3.52 1.22 3.575 1.56 ;
      RECT 3.52 3.135 3.575 3.945 ;
      RECT 3.1 1.325 3.14 1.665 ;
      RECT 2.87 0.63 3.1 1.095 ;
      RECT 2.87 1.325 3.1 4.405 ;
      RECT 0.52 0.865 2.87 1.095 ;
      RECT 2.8 1.325 2.87 1.665 ;
      RECT 2.76 2.74 2.87 3.08 ;
      RECT 1.84 2.04 2.585 2.38 ;
      RECT 1.61 1.46 1.84 3.08 ;
      RECT 1.5 1.46 1.61 1.8 ;
      RECT 1.5 2.74 1.61 3.08 ;
      RECT 0.29 0.865 0.52 3.08 ;
      RECT 0.18 1.46 0.29 1.8 ;
      RECT 0.18 2.74 0.29 3.08 ;
  END
END AFCSHCONX2

MACRO AFCSHCINX4
  CLASS CORE ;
  FOREIGN AFCSHCINX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 32.34 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 1.1475 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1552 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 32.2 0.97 32.21 3.025 ;
      RECT 31.98 0.97 32.2 4.34 ;
      RECT 31.82 0.97 31.98 1.78 ;
      RECT 31.82 2.74 31.98 4.34 ;
     END
  END S

  PIN CS
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.44 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0935 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 31.13 1.26 31.54 1.54 ;
      RECT 30.9 1.26 31.13 2.43 ;
      RECT 30.735 2.09 30.9 2.43 ;
     END
  END CS

  PIN CO1
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.522 ;
  ANTENNAPARTIALMETALAREA 2.1685 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.3386 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 18.34 2.205 21.7 2.435 ;
      RECT 18.34 3.685 21.7 3.915 ;
      RECT 18.055 2.205 18.34 3.915 ;
      RECT 18.035 2.38 18.055 3.915 ;
      RECT 17.96 2.38 18.035 3.78 ;
     END
  END CO1

  PIN CO0
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.513 ;
  ANTENNAPARTIALMETALAREA 2.1583 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.2326 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.635 2.38 17.68 3.78 ;
      RECT 17.3 2.205 17.635 3.915 ;
      RECT 13.99 2.205 17.3 2.435 ;
      RECT 13.99 3.685 17.3 3.915 ;
     END
  END CO0

  PIN CI1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0194 ;
  ANTENNAPARTIALMETALAREA 0.2227 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0017 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 25.88 2.28 26.375 2.73 ;
     END
  END CI1N

  PIN CI0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9978 ;
  ANTENNAPARTIALMETALAREA 0.207 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9699 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.38 2.25 9.885 2.66 ;
     END
  END CI0N

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5034 ;
  ANTENNAPARTIALMETALAREA 0.2291 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.715 2.315 9.1 2.91 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.759 ;
  ANTENNAPARTIALMETALAREA 0.2881 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5158 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.105 1.18 2.445 ;
      RECT 0.875 2.105 1.105 3.195 ;
      RECT 0.84 2.105 0.875 2.445 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 31.4 -0.4 32.34 0.4 ;
      RECT 31.06 -0.4 31.4 0.63 ;
      RECT 29.87 -0.4 31.06 0.4 ;
      RECT 29.53 -0.4 29.87 1.78 ;
      RECT 26.695 -0.4 29.53 0.4 ;
      RECT 26.355 -0.4 26.695 0.575 ;
      RECT 25.335 -0.4 26.355 0.4 ;
      RECT 24.995 -0.4 25.335 0.575 ;
      RECT 10.725 -0.4 24.995 0.4 ;
      RECT 10.385 -0.4 10.725 0.575 ;
      RECT 9.335 -0.4 10.385 0.4 ;
      RECT 8.995 -0.4 9.335 0.575 ;
      RECT 7.945 -0.4 8.995 0.4 ;
      RECT 7.605 -0.4 7.945 0.575 ;
      RECT 2.38 -0.4 7.605 0.4 ;
      RECT 2.04 -0.4 2.38 0.63 ;
      RECT 1.2 -0.4 2.04 0.4 ;
      RECT 0.86 -0.4 1.2 0.63 ;
      RECT 0 -0.4 0.86 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 31.48 4.64 32.34 5.44 ;
      RECT 31.14 3.94 31.48 5.44 ;
      RECT 30.535 4.64 31.14 5.44 ;
      RECT 30.195 3.76 30.535 5.44 ;
      RECT 26.695 4.64 30.195 5.44 ;
      RECT 26.355 4.465 26.695 5.44 ;
      RECT 25.335 4.64 26.355 5.44 ;
      RECT 24.995 4.465 25.335 5.44 ;
      RECT 10.725 4.64 24.995 5.44 ;
      RECT 10.385 4.465 10.725 5.44 ;
      RECT 9.335 4.64 10.385 5.44 ;
      RECT 8.995 4.465 9.335 5.44 ;
      RECT 7.945 4.64 8.995 5.44 ;
      RECT 7.605 4.465 7.945 5.44 ;
      RECT 2.38 4.64 7.605 5.44 ;
      RECT 2.04 3.94 2.38 5.44 ;
      RECT 1.16 4.64 2.04 5.44 ;
      RECT 0.82 4.09 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 31.59 2.17 31.75 2.51 ;
      RECT 31.36 2.17 31.59 3.505 ;
      RECT 29.96 3.275 31.36 3.505 ;
      RECT 30.5 1.46 30.665 1.8 ;
      RECT 30.5 2.795 30.665 3.025 ;
      RECT 30.27 1.46 30.5 3.025 ;
      RECT 29.5 2.795 30.27 3.025 ;
      RECT 29.73 3.275 29.96 4.405 ;
      RECT 28.12 4.175 29.73 4.405 ;
      RECT 29.27 2.795 29.5 3.915 ;
      RECT 29.3 2.095 29.41 2.325 ;
      RECT 29.07 0.815 29.3 2.325 ;
      RECT 28.58 3.685 29.27 3.915 ;
      RECT 22.495 0.815 29.07 1.045 ;
      RECT 28.84 2.62 29.04 3.445 ;
      RECT 28.81 1.38 28.84 3.445 ;
      RECT 28.61 1.38 28.81 2.85 ;
      RECT 28.38 3.08 28.58 3.915 ;
      RECT 28.35 2.17 28.38 3.915 ;
      RECT 28.15 2.17 28.35 3.31 ;
      RECT 27.915 1.38 28.175 1.72 ;
      RECT 27.915 3.54 28.12 4.405 ;
      RECT 27.89 1.38 27.915 4.405 ;
      RECT 27.685 1.38 27.89 3.77 ;
      RECT 27.225 1.38 27.455 3.965 ;
      RECT 27.115 1.38 27.225 1.72 ;
      RECT 27.115 3.155 27.225 3.965 ;
      RECT 26.835 2.39 26.945 2.73 ;
      RECT 26.605 1.275 26.835 2.73 ;
      RECT 23.96 1.275 26.605 1.505 ;
      RECT 25.645 1.735 26.015 1.965 ;
      RECT 25.64 2.96 25.96 3.775 ;
      RECT 25.64 1.735 25.645 2.665 ;
      RECT 25.41 1.735 25.64 3.775 ;
      RECT 24.715 2.435 25.41 2.665 ;
      RECT 22.955 3.545 25.41 3.775 ;
      RECT 24.445 3.08 24.625 3.31 ;
      RECT 24.445 1.735 24.615 1.965 ;
      RECT 24.215 1.735 24.445 3.31 ;
      RECT 11.59 4.18 24.385 4.41 ;
      RECT 23.73 1.275 23.96 3.25 ;
      RECT 23.515 1.275 23.73 1.505 ;
      RECT 23.565 3.02 23.73 3.25 ;
      RECT 22.955 1.385 23.08 1.615 ;
      RECT 22.725 1.385 22.955 3.775 ;
      RECT 18.75 2.965 22.725 3.195 ;
      RECT 22.265 0.815 22.495 1.965 ;
      RECT 13.24 1.735 22.265 1.965 ;
      RECT 20.09 0.74 22.03 0.97 ;
      RECT 7.185 1.265 21.7 1.495 ;
      RECT 19.805 0.735 20.09 0.97 ;
      RECT 11.21 0.735 19.805 0.965 ;
      RECT 13.295 2.965 16.94 3.195 ;
      RECT 13.295 2.195 13.405 2.425 ;
      RECT 13.065 2.195 13.295 3.79 ;
      RECT 13.01 1.725 13.24 1.965 ;
      RECT 12.83 3.56 13.065 3.79 ;
      RECT 12.16 1.725 13.01 1.955 ;
      RECT 12.545 3.545 12.83 3.79 ;
      RECT 10.265 3.545 12.545 3.775 ;
      RECT 11.93 1.725 12.16 3.31 ;
      RECT 11.835 1.725 11.93 1.955 ;
      RECT 11.785 3.08 11.93 3.31 ;
      RECT 11.305 4.005 11.59 4.41 ;
      RECT 11.245 1.725 11.475 3.31 ;
      RECT 4.65 4.005 11.305 4.235 ;
      RECT 11.115 1.725 11.245 1.955 ;
      RECT 11.065 3.08 11.245 3.31 ;
      RECT 10.98 0.735 11.21 1.035 ;
      RECT 7.28 0.805 10.98 1.035 ;
      RECT 10.535 2.435 10.975 2.665 ;
      RECT 10.305 1.725 10.535 3.18 ;
      RECT 9.705 1.725 10.305 1.955 ;
      RECT 10.265 2.95 10.305 3.18 ;
      RECT 9.76 2.95 10.265 3.775 ;
      RECT 8.46 1.725 8.655 1.955 ;
      RECT 8.46 3.165 8.655 3.505 ;
      RECT 8.315 1.725 8.46 3.505 ;
      RECT 8.23 1.725 8.315 3.45 ;
      RECT 7.405 2.185 8.23 2.54 ;
      RECT 7.05 0.63 7.28 1.035 ;
      RECT 7.075 1.265 7.185 1.825 ;
      RECT 7.075 2.955 7.185 3.295 ;
      RECT 6.845 1.265 7.075 3.295 ;
      RECT 5.245 0.63 7.05 0.86 ;
      RECT 6.575 1.265 6.845 1.495 ;
      RECT 6.59 3.065 6.845 3.295 ;
      RECT 6.36 3.065 6.59 3.76 ;
      RECT 6.235 1.12 6.575 1.495 ;
      RECT 6.25 3.42 6.36 3.76 ;
      RECT 5.775 1.205 6.005 3.575 ;
      RECT 5.735 1.205 5.775 1.665 ;
      RECT 3.14 3.345 5.775 3.575 ;
      RECT 5.245 2.765 5.34 3.105 ;
      RECT 5.015 0.63 5.245 3.105 ;
      RECT 5 2.765 5.015 3.105 ;
      RECT 4.42 3.81 4.65 4.235 ;
      RECT 4.51 2.765 4.62 3.105 ;
      RECT 4.51 1.075 4.58 1.415 ;
      RECT 4.47 1.075 4.51 3.105 ;
      RECT 4.28 0.63 4.47 3.105 ;
      RECT 3.56 3.81 4.42 4.04 ;
      RECT 4.24 0.63 4.28 1.415 ;
      RECT 3.1 0.63 4.24 0.86 ;
      RECT 3.79 2.76 3.9 3.1 ;
      RECT 3.79 1.22 3.86 1.56 ;
      RECT 3.56 1.22 3.79 3.1 ;
      RECT 3.52 1.22 3.56 1.56 ;
      RECT 2.91 1.325 3.14 4.015 ;
      RECT 2.87 0.63 3.1 1.095 ;
      RECT 2.8 1.325 2.91 1.665 ;
      RECT 2.8 3.205 2.91 4.015 ;
      RECT 0.52 0.865 2.87 1.095 ;
      RECT 1.84 2.04 2.585 2.38 ;
      RECT 1.61 1.46 1.84 3.395 ;
      RECT 1.5 1.46 1.61 1.8 ;
      RECT 1.5 3.055 1.61 3.395 ;
      RECT 0.29 0.865 0.52 3.08 ;
      RECT 0.18 1.46 0.29 1.8 ;
      RECT 0.18 2.74 0.29 3.08 ;
  END
END AFCSHCINX4

MACRO AFCSHCINX2
  CLASS CORE ;
  FOREIGN AFCSHCINX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 29.7 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AFCSHCINX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3356 ;
  ANTENNAPARTIALMETALAREA 1.1475 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1552 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 29.56 0.97 29.57 3.025 ;
      RECT 29.34 0.97 29.56 4.34 ;
      RECT 29.18 0.97 29.34 1.78 ;
      RECT 29.18 2.74 29.34 4.34 ;
     END
  END S

  PIN CS
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5814 ;
  ANTENNAPARTIALMETALAREA 0.44 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0935 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 28.49 1.26 28.9 1.54 ;
      RECT 28.26 1.26 28.49 2.43 ;
      RECT 28.095 2.09 28.26 2.43 ;
     END
  END CS

  PIN CO1
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.3194 ;
  ANTENNAPARTIALMETALAREA 1.1931 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.3212 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 19 3.48 19.735 3.71 ;
      RECT 19 2.2 19.515 2.43 ;
      RECT 18.77 2.2 19 3.78 ;
      RECT 18.62 2.94 18.77 3.78 ;
      RECT 17.62 3.48 18.62 3.71 ;
      RECT 17.39 3.135 17.62 3.945 ;
     END
  END CO1

  PIN CO0
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.3194 ;
  ANTENNAPARTIALMETALAREA 1.1437 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.0933 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.55 3.135 15.78 3.945 ;
      RECT 14.38 3.48 15.55 3.71 ;
      RECT 14.23 2.94 14.38 3.78 ;
      RECT 14 2.195 14.23 3.78 ;
      RECT 13.655 2.195 14 2.425 ;
      RECT 13.485 3.48 14 3.71 ;
     END
  END CO0

  PIN CI1N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5097 ;
  ANTENNAPARTIALMETALAREA 0.2295 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 23.735 2.39 23.755 2.73 ;
      RECT 23.24 2.28 23.735 2.73 ;
     END
  END CI1N

  PIN CI0N
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5079 ;
  ANTENNAPARTIALMETALAREA 0.2284 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0176 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.38 2.195 9.815 2.72 ;
     END
  END CI0N

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5034 ;
  ANTENNAPARTIALMETALAREA 0.2328 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.615 2.22 9.1 2.7 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7626 ;
  ANTENNAPARTIALMETALAREA 0.2881 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.5158 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.105 2.105 1.18 2.445 ;
      RECT 0.875 2.105 1.105 3.195 ;
      RECT 0.84 2.105 0.875 2.445 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 28.76 -0.4 29.7 0.4 ;
      RECT 28.42 -0.4 28.76 0.63 ;
      RECT 27.24 -0.4 28.42 0.4 ;
      RECT 27.01 -0.4 27.24 1.78 ;
      RECT 24.175 -0.4 27.01 0.4 ;
      RECT 23.835 -0.4 24.175 0.575 ;
      RECT 22.745 -0.4 23.835 0.4 ;
      RECT 22.405 -0.4 22.745 0.575 ;
      RECT 10.765 -0.4 22.405 0.4 ;
      RECT 10.425 -0.4 10.765 0.575 ;
      RECT 9.305 -0.4 10.425 0.4 ;
      RECT 8.965 -0.4 9.305 0.575 ;
      RECT 7.925 -0.4 8.965 0.4 ;
      RECT 7.585 -0.4 7.925 0.575 ;
      RECT 2.35 -0.4 7.585 0.4 ;
      RECT 2.01 -0.4 2.35 0.63 ;
      RECT 1.17 -0.4 2.01 0.4 ;
      RECT 0.83 -0.4 1.17 0.63 ;
      RECT 0 -0.4 0.83 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 28.84 4.64 29.7 5.44 ;
      RECT 28.5 3.94 28.84 5.44 ;
      RECT 28.015 4.64 28.5 5.44 ;
      RECT 27.675 3.76 28.015 5.44 ;
      RECT 24.175 4.64 27.675 5.44 ;
      RECT 23.835 4.465 24.175 5.44 ;
      RECT 22.795 4.64 23.835 5.44 ;
      RECT 22.455 4.465 22.795 5.44 ;
      RECT 10.715 4.64 22.455 5.44 ;
      RECT 10.375 4.465 10.715 5.44 ;
      RECT 9.305 4.64 10.375 5.44 ;
      RECT 8.965 4.465 9.305 5.44 ;
      RECT 7.925 4.64 8.965 5.44 ;
      RECT 7.585 4.465 7.925 5.44 ;
      RECT 2.39 4.64 7.585 5.44 ;
      RECT 2.05 3.94 2.39 5.44 ;
      RECT 1.16 4.64 2.05 5.44 ;
      RECT 0.82 3.81 1.16 5.44 ;
      RECT 0 4.64 0.82 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 28.95 2.17 29.11 2.51 ;
      RECT 28.72 2.17 28.95 3.505 ;
      RECT 27.44 3.275 28.72 3.505 ;
      RECT 27.85 1.46 28.015 1.8 ;
      RECT 27.85 2.795 28.015 3.025 ;
      RECT 27.62 1.46 27.85 3.025 ;
      RECT 26.98 2.795 27.62 3.025 ;
      RECT 27.21 3.275 27.44 4.405 ;
      RECT 25.6 4.175 27.21 4.405 ;
      RECT 26.75 2.795 26.98 3.915 ;
      RECT 26.78 2.095 26.89 2.325 ;
      RECT 26.55 0.815 26.78 2.325 ;
      RECT 26.06 3.685 26.75 3.915 ;
      RECT 20.99 0.815 26.55 1.045 ;
      RECT 26.32 2.62 26.52 3.45 ;
      RECT 26.29 1.38 26.32 3.45 ;
      RECT 26.09 1.38 26.29 2.85 ;
      RECT 25.86 3.08 26.06 3.915 ;
      RECT 25.83 2.17 25.86 3.915 ;
      RECT 25.63 2.17 25.83 3.31 ;
      RECT 25.395 1.38 25.655 1.72 ;
      RECT 25.395 3.54 25.6 4.405 ;
      RECT 25.37 1.38 25.395 4.405 ;
      RECT 25.165 1.38 25.37 3.77 ;
      RECT 24.705 1.38 24.935 3.965 ;
      RECT 24.595 1.38 24.705 1.72 ;
      RECT 24.595 3.155 24.705 3.965 ;
      RECT 24.315 2.39 24.425 2.73 ;
      RECT 24.085 1.275 24.315 2.73 ;
      RECT 21.515 1.275 24.085 1.505 ;
      RECT 23.01 1.735 23.495 1.965 ;
      RECT 23.01 2.96 23.44 3.8 ;
      RECT 22.78 1.735 23.01 3.8 ;
      RECT 22.325 2.435 22.78 2.665 ;
      RECT 20.7 3.57 22.78 3.8 ;
      RECT 22.055 3.08 22.235 3.31 ;
      RECT 22.055 1.735 22.185 1.965 ;
      RECT 21.825 1.735 22.055 3.31 ;
      RECT 11.23 4.18 21.995 4.41 ;
      RECT 21.285 1.275 21.515 3.31 ;
      RECT 20.655 1.735 21.285 1.965 ;
      RECT 21.175 3.08 21.285 3.31 ;
      RECT 20.76 0.815 20.99 1.485 ;
      RECT 19.455 1.255 20.76 1.485 ;
      RECT 20.47 2.2 20.7 3.8 ;
      RECT 19.895 2.2 20.47 2.43 ;
      RECT 19.82 0.74 19.875 0.97 ;
      RECT 19.59 0.735 19.82 0.97 ;
      RECT 11.265 0.735 19.59 0.965 ;
      RECT 19.225 1.255 19.455 1.965 ;
      RECT 17.16 1.735 19.225 1.965 ;
      RECT 18.7 1.275 18.755 1.505 ;
      RECT 16.7 1.265 18.7 1.505 ;
      RECT 16.93 1.735 17.16 3.5 ;
      RECT 16.24 3.27 16.93 3.5 ;
      RECT 16.47 1.265 16.7 3.035 ;
      RECT 7.165 1.265 16.47 1.495 ;
      RECT 16.01 1.775 16.24 3.5 ;
      RECT 14.855 1.775 16.01 2.005 ;
      RECT 14.625 1.735 14.855 2.005 ;
      RECT 12.03 1.735 14.625 1.965 ;
      RECT 12.7 2.195 13.275 2.425 ;
      RECT 12.47 2.195 12.7 3.775 ;
      RECT 10.32 3.545 12.47 3.775 ;
      RECT 11.8 1.735 12.03 3.31 ;
      RECT 11.705 1.735 11.8 1.965 ;
      RECT 11.655 3.08 11.8 3.31 ;
      RECT 11.115 1.735 11.345 3.31 ;
      RECT 11.035 0.735 11.265 1.035 ;
      RECT 11 4.005 11.23 4.41 ;
      RECT 10.985 1.735 11.115 1.965 ;
      RECT 10.935 3.08 11.115 3.31 ;
      RECT 7.29 0.805 11.035 1.035 ;
      RECT 3.885 4.005 11 4.235 ;
      RECT 10.32 2.435 10.845 2.665 ;
      RECT 10.09 1.735 10.32 3.775 ;
      RECT 9.675 1.735 10.09 1.965 ;
      RECT 9.73 2.95 10.09 3.775 ;
      RECT 8.385 1.73 8.625 1.96 ;
      RECT 8.385 2.95 8.57 3.775 ;
      RECT 8.34 1.73 8.385 3.775 ;
      RECT 8.155 1.73 8.34 3.18 ;
      RECT 7.385 2.185 8.155 2.525 ;
      RECT 7.06 0.63 7.29 1.035 ;
      RECT 7.11 1.265 7.165 1.605 ;
      RECT 6.88 1.265 7.11 3.765 ;
      RECT 5.255 0.63 7.06 0.86 ;
      RECT 6.825 1.265 6.88 1.605 ;
      RECT 6.245 3.42 6.88 3.765 ;
      RECT 6.585 1.265 6.825 1.495 ;
      RECT 6.245 1.12 6.585 1.495 ;
      RECT 5.745 1.235 5.975 3.6 ;
      RECT 3.07 3.365 5.745 3.595 ;
      RECT 5.025 0.63 5.255 3.135 ;
      RECT 4.48 1.075 4.59 1.415 ;
      RECT 4.48 2.795 4.59 3.135 ;
      RECT 4.44 1.075 4.48 3.135 ;
      RECT 4.25 0.63 4.44 3.135 ;
      RECT 4.21 0.63 4.25 1.36 ;
      RECT 3.1 0.63 4.21 0.86 ;
      RECT 3.53 3.825 3.885 4.235 ;
      RECT 3.815 1.22 3.87 1.56 ;
      RECT 3.815 2.795 3.87 3.135 ;
      RECT 3.585 1.22 3.815 3.135 ;
      RECT 3.53 1.22 3.585 1.56 ;
      RECT 3.53 2.795 3.585 3.135 ;
      RECT 3.07 1.325 3.15 1.665 ;
      RECT 2.87 0.63 3.1 1.095 ;
      RECT 2.84 1.325 3.07 3.595 ;
      RECT 0.52 0.865 2.87 1.095 ;
      RECT 2.81 1.325 2.84 1.665 ;
      RECT 2.73 2.85 2.84 3.19 ;
      RECT 1.78 2.04 2.555 2.38 ;
      RECT 1.78 1.46 1.84 1.8 ;
      RECT 1.78 2.74 1.81 3.08 ;
      RECT 1.55 1.46 1.78 3.08 ;
      RECT 1.5 1.46 1.55 1.8 ;
      RECT 1.47 2.74 1.55 3.08 ;
      RECT 0.29 0.865 0.52 3.08 ;
      RECT 0.18 1.46 0.29 1.8 ;
      RECT 0.18 2.74 0.29 3.08 ;
  END
END AFCSHCINX2

MACRO AHHCONX4
  CLASS CORE ;
  FOREIGN AHHCONX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.58 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.0254 ;
  ANTENNAPARTIALMETALAREA 1.1292 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.5792 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.33 1.82 4.48 3.22 ;
      RECT 4.1 1.33 4.33 3.22 ;
      RECT 3.935 1.33 4.1 1.56 ;
      RECT 3.515 2.84 4.1 3.07 ;
      RECT 3.615 1.21 3.935 1.56 ;
      RECT 3.5 2.84 3.515 3.22 ;
      RECT 3.27 2.84 3.5 3.685 ;
     END
  END S

  PIN CON
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.2774 ;
  ANTENNAPARTIALMETALAREA 2.5319 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.6549 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.42 1.82 8.44 3.22 ;
      RECT 8.06 1.365 8.42 3.43 ;
      RECT 6.815 1.365 8.06 1.595 ;
      RECT 7.445 3.09 8.06 3.43 ;
      RECT 7.105 3.09 7.445 3.9 ;
      RECT 5.96 3.09 7.105 3.43 ;
      RECT 6.7 1.26 6.815 1.595 ;
      RECT 6.36 0.705 6.7 1.595 ;
      RECT 5.64 3.09 5.96 3.9 ;
     END
  END CON

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.6038 ;
  ANTENNAPARTIALMETALAREA 2.4702 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.5152 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.095 2.29 6.94 2.69 ;
      RECT 5.41 2.46 6.095 2.69 ;
      RECT 5.18 2.46 5.41 4.145 ;
      RECT 3.04 3.915 5.18 4.145 ;
      RECT 3.64 1.8 3.87 2.52 ;
      RECT 3.04 2.29 3.64 2.52 ;
      RECT 2.81 2.29 3.04 4.145 ;
      RECT 2.215 2.29 2.81 2.66 ;
      RECT 1.875 2.235 2.215 2.66 ;
     END
  END CI

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3932 ;
  ANTENNAPARTIALMETALAREA 0.7849 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6888 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.345 1.83 7.685 2.23 ;
      RECT 5.725 1.83 7.345 2.06 ;
      RECT 5.66 1.285 5.725 2.06 ;
      RECT 5.495 1.285 5.66 2.23 ;
      RECT 5.32 1.83 5.495 2.23 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.02 -0.4 8.58 0.4 ;
      RECT 7.68 -0.4 8.02 1.105 ;
      RECT 5.38 -0.4 7.68 0.4 ;
      RECT 5.04 -0.4 5.38 0.575 ;
      RECT 1.34 -0.4 5.04 0.4 ;
      RECT 1 -0.4 1.34 0.575 ;
      RECT 0 -0.4 1 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 8.245 4.64 8.58 5.44 ;
      RECT 7.905 3.935 8.245 5.44 ;
      RECT 6.685 4.64 7.905 5.44 ;
      RECT 6.345 3.935 6.685 5.44 ;
      RECT 5.035 4.64 6.345 5.44 ;
      RECT 4.695 4.41 5.035 5.44 ;
      RECT 1.335 4.64 4.695 5.44 ;
      RECT 0.995 4.41 1.335 5.44 ;
      RECT 0 4.64 0.995 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 4.72 0.81 4.95 3.685 ;
      RECT 4.62 0.81 4.72 1.04 ;
      RECT 3.935 3.455 4.72 3.685 ;
      RECT 4.28 0.675 4.62 1.04 ;
      RECT 3.385 0.73 4.28 0.96 ;
      RECT 3.155 0.73 3.385 1.955 ;
      RECT 1.49 1.725 3.155 1.955 ;
      RECT 2.6 0.63 2.925 1.035 ;
      RECT 1.03 1.265 2.68 1.495 ;
      RECT 0.57 0.805 2.6 1.035 ;
      RECT 2.215 3.92 2.53 4.29 ;
      RECT 0.57 3.92 2.215 4.15 ;
      RECT 1.705 3.18 2.045 3.52 ;
      RECT 1.03 3.18 1.705 3.41 ;
      RECT 1.26 1.725 1.49 2.56 ;
      RECT 0.8 1.265 1.03 3.41 ;
      RECT 0.23 0.76 0.57 4.15 ;
  END
END AHHCONX4

MACRO AHHCONX2
  CLASS CORE ;
  FOREIGN AHHCONX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AHHCONX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.7726 ;
  ANTENNAPARTIALMETALAREA 1.0937 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.6004 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.26 1.33 4.49 3.22 ;
      RECT 3.845 1.33 4.26 1.56 ;
      RECT 3.5 2.84 4.26 3.22 ;
      RECT 3.615 1.21 3.845 1.56 ;
      RECT 3.27 2.84 3.5 3.685 ;
     END
  END S

  PIN CON
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4296 ;
  ANTENNAPARTIALMETALAREA 1.3379 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.5067 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.815 1.285 7.045 4.04 ;
      RECT 6.7 1.26 6.815 1.515 ;
      RECT 5.64 3.7 6.815 4.04 ;
      RECT 6.36 0.705 6.7 1.515 ;
     END
  END CON

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.1322 ;
  ANTENNAPARTIALMETALAREA 2.2151 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.9216 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.09 2.235 6.32 3.3 ;
      RECT 5.41 3.07 6.09 3.3 ;
      RECT 5.18 3.07 5.41 4.145 ;
      RECT 3.04 3.915 5.18 4.145 ;
      RECT 3.8 1.8 4.03 2.52 ;
      RECT 3.04 2.29 3.8 2.52 ;
      RECT 2.81 2.29 3.04 4.145 ;
      RECT 2.37 2.29 2.81 2.66 ;
      RECT 2.03 2.235 2.37 2.66 ;
     END
  END CI

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9216 ;
  ANTENNAPARTIALMETALAREA 0.3107 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1819 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.76 1.74 5.315 2.3 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.38 -0.4 7.26 0.4 ;
      RECT 5.04 -0.4 5.38 0.575 ;
      RECT 1.34 -0.4 5.04 0.4 ;
      RECT 1 -0.4 1.34 0.575 ;
      RECT 0 -0.4 1 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.685 4.64 7.26 5.44 ;
      RECT 6.345 4.41 6.685 5.44 ;
      RECT 5.035 4.64 6.345 5.44 ;
      RECT 4.695 4.41 5.035 5.44 ;
      RECT 1.335 4.64 4.695 5.44 ;
      RECT 0.995 4.41 1.335 5.44 ;
      RECT 0 4.64 0.995 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.565 0.81 5.795 2.825 ;
      RECT 4.62 0.81 5.565 1.04 ;
      RECT 4.95 2.595 5.565 2.825 ;
      RECT 4.72 2.595 4.95 3.685 ;
      RECT 3.935 3.455 4.72 3.685 ;
      RECT 4.28 0.675 4.62 1.04 ;
      RECT 3.385 0.73 4.28 0.96 ;
      RECT 3.155 0.73 3.385 1.955 ;
      RECT 1.605 1.725 3.155 1.955 ;
      RECT 2.6 0.63 2.925 1.035 ;
      RECT 1.035 1.265 2.805 1.495 ;
      RECT 0.575 0.805 2.6 1.035 ;
      RECT 2.265 3.92 2.58 4.29 ;
      RECT 0.575 3.92 2.265 4.15 ;
      RECT 1.755 3.18 2.095 3.52 ;
      RECT 1.035 3.18 1.755 3.41 ;
      RECT 1.375 1.725 1.605 2.56 ;
      RECT 1.265 2.22 1.375 2.56 ;
      RECT 0.805 1.265 1.035 3.41 ;
      RECT 0.235 0.76 0.575 4.15 ;
  END
END AHHCONX2

MACRO AHHCINX4
  CLASS CORE ;
  FOREIGN AHHCINX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.92 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5924 ;
  ANTENNAPARTIALMETALAREA 1.0118 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.6941 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.215 2.91 3.555 3.73 ;
      RECT 3.18 1.27 3.41 2.05 ;
      RECT 3.16 2.91 3.215 3.22 ;
      RECT 3.16 1.82 3.18 2.05 ;
      RECT 2.78 1.82 3.16 3.22 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.8914 ;
  ANTENNAPARTIALMETALAREA 1.7415 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.3653 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.02 1.82 7.12 3.22 ;
      RECT 6.74 0.99 7.02 3.22 ;
      RECT 6.68 0.99 6.74 1.8 ;
      RECT 6.42 2.78 6.74 3.01 ;
      RECT 6.385 1.26 6.68 1.56 ;
      RECT 6.08 2.78 6.42 3.59 ;
      RECT 5.625 1.33 6.385 1.56 ;
      RECT 5.285 0.63 5.625 1.56 ;
     END
  END CO

  PIN CIN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.5858 ;
  ANTENNAPARTIALMETALAREA 2.336 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.9498 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.58 2.13 7.69 2.47 ;
      RECT 7.35 2.13 7.58 3.68 ;
      RECT 6.88 3.45 7.35 3.68 ;
      RECT 6.65 3.45 6.88 4.05 ;
      RECT 5.8 3.82 6.65 4.05 ;
      RECT 5.785 3.78 5.8 4.05 ;
      RECT 5.555 3.48 5.785 4.05 ;
      RECT 5.295 3.48 5.555 3.71 ;
      RECT 5.065 2.25 5.295 3.71 ;
      RECT 4.41 3.48 5.065 3.71 ;
      RECT 4.18 3.48 4.41 4.37 ;
      RECT 4.175 4.085 4.18 4.37 ;
      RECT 1.51 4.14 4.175 4.37 ;
     END
  END CIN

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4338 ;
  ANTENNAPARTIALMETALAREA 0.349 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.265 1.8 4.375 2.14 ;
      RECT 4.035 1.8 4.265 2.61 ;
      RECT 3.745 2.38 4.035 2.61 ;
      RECT 3.515 2.38 3.745 2.635 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.74 -0.4 7.92 0.4 ;
      RECT 7.4 -0.4 7.74 1.8 ;
      RECT 6.385 -0.4 7.4 0.4 ;
      RECT 6.045 -0.4 6.385 0.63 ;
      RECT 4.905 -0.4 6.045 0.4 ;
      RECT 4.565 -0.4 4.905 0.97 ;
      RECT 1.28 -0.4 4.565 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.74 4.64 7.92 5.44 ;
      RECT 7.4 3.94 7.74 5.44 ;
      RECT 5.05 4.64 7.4 5.44 ;
      RECT 4.71 3.94 5.05 5.44 ;
      RECT 1.28 4.64 4.71 5.44 ;
      RECT 0.94 4.41 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.91 1.99 6.02 2.33 ;
      RECT 5.68 1.79 5.91 2.33 ;
      RECT 4.835 1.79 5.68 2.02 ;
      RECT 4.605 1.28 4.835 3.25 ;
      RECT 4.185 1.28 4.605 1.51 ;
      RECT 3.935 2.91 4.605 3.25 ;
      RECT 3.845 0.7 4.185 1.51 ;
      RECT 2.95 0.75 3.845 0.98 ;
      RECT 2.72 0.75 2.95 1.495 ;
      RECT 2.455 3.57 2.795 3.91 ;
      RECT 2.405 1.265 2.72 1.495 ;
      RECT 2.18 0.63 2.49 1.035 ;
      RECT 0.52 3.68 2.455 3.91 ;
      RECT 2.085 2.23 2.425 2.57 ;
      RECT 2.175 1.265 2.405 1.955 ;
      RECT 0.52 0.805 2.18 1.035 ;
      RECT 1.27 1.725 2.175 1.955 ;
      RECT 1.88 2.34 2.085 2.57 ;
      RECT 1.65 2.34 1.88 3.45 ;
      RECT 0.81 1.265 1.845 1.495 ;
      RECT 1.54 3.11 1.65 3.45 ;
      RECT 0.81 3.11 1.54 3.34 ;
      RECT 1.04 1.725 1.27 2.5 ;
      RECT 0.58 1.265 0.81 3.34 ;
      RECT 0.35 0.695 0.52 1.035 ;
      RECT 0.35 3.61 0.52 3.95 ;
      RECT 0.12 0.695 0.35 3.95 ;
  END
END AHHCINX4

MACRO AHHCINX2
  CLASS CORE ;
  FOREIGN AHHCINX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AHHCINX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.5924 ;
  ANTENNAPARTIALMETALAREA 0.853 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7471 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.215 2.91 3.555 3.73 ;
      RECT 3.18 1.21 3.41 1.955 ;
      RECT 3.095 2.91 3.215 3.22 ;
      RECT 3.095 1.725 3.18 1.955 ;
      RECT 2.865 1.725 3.095 3.22 ;
      RECT 2.855 2.405 2.865 2.635 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.254 ;
  ANTENNAPARTIALMETALAREA 1.2814 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.0456 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.42 1.33 6.48 2.66 ;
      RECT 6.25 1.33 6.42 4.06 ;
      RECT 5.66 1.33 6.25 1.56 ;
      RECT 6.08 2.38 6.25 4.06 ;
      RECT 5.32 0.63 5.66 1.56 ;
     END
  END CO

  PIN CIN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.143 ;
  ANTENNAPARTIALMETALAREA 1.3055 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.2593 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.065 2.25 5.295 3.71 ;
      RECT 4.41 3.48 5.065 3.71 ;
      RECT 4.18 3.48 4.41 4.37 ;
      RECT 4.175 4.085 4.18 4.37 ;
      RECT 1.51 4.14 4.175 4.37 ;
     END
  END CIN

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4338 ;
  ANTENNAPARTIALMETALAREA 0.349 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.7967 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.265 1.8 4.375 2.14 ;
      RECT 4.035 1.8 4.265 2.61 ;
      RECT 3.745 2.38 4.035 2.61 ;
      RECT 3.515 2.38 3.745 2.635 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.42 -0.4 6.6 0.4 ;
      RECT 6.08 -0.4 6.42 1.1 ;
      RECT 4.905 -0.4 6.08 0.4 ;
      RECT 4.565 -0.4 4.905 0.97 ;
      RECT 1.285 -0.4 4.565 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 5.05 4.64 6.6 5.44 ;
      RECT 4.71 3.94 5.05 5.44 ;
      RECT 1.28 4.64 4.71 5.44 ;
      RECT 0.94 4.41 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 5.68 1.79 6.02 2.13 ;
      RECT 4.835 1.79 5.68 2.02 ;
      RECT 4.605 1.28 4.835 3.25 ;
      RECT 4.185 1.28 4.605 1.51 ;
      RECT 3.935 2.91 4.605 3.25 ;
      RECT 3.845 0.7 4.185 1.51 ;
      RECT 2.95 0.75 3.845 0.98 ;
      RECT 2.72 0.75 2.95 1.495 ;
      RECT 2.405 1.265 2.72 1.495 ;
      RECT 2.295 3.1 2.635 3.91 ;
      RECT 2.165 0.63 2.49 1.035 ;
      RECT 2.085 2.23 2.425 2.57 ;
      RECT 2.175 1.265 2.405 1.955 ;
      RECT 0.52 3.68 2.295 3.91 ;
      RECT 1.27 1.725 2.175 1.955 ;
      RECT 0.52 0.805 2.165 1.035 ;
      RECT 1.88 2.34 2.085 2.57 ;
      RECT 1.65 2.34 1.88 3.45 ;
      RECT 0.81 1.265 1.845 1.495 ;
      RECT 1.54 3.11 1.65 3.45 ;
      RECT 0.81 3.11 1.54 3.34 ;
      RECT 1.04 1.725 1.27 2.5 ;
      RECT 0.58 1.265 0.81 3.34 ;
      RECT 0.35 0.695 0.52 1.035 ;
      RECT 0.35 3.61 0.52 3.95 ;
      RECT 0.12 0.695 0.35 3.95 ;
  END
END AHHCINX2

MACRO AFHCONX4
  CLASS CORE ;
  FOREIGN AFHCONX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1328 ;
  ANTENNAPARTIALMETALAREA 1.1633 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.4255 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.58 1.82 15.7 3.22 ;
      RECT 15.32 1.515 15.58 3.22 ;
      RECT 15.3 1.515 15.32 1.775 ;
      RECT 14.985 2.815 15.32 3.045 ;
      RECT 14.96 0.965 15.3 1.775 ;
      RECT 14.755 2.815 14.985 3.66 ;
     END
  END S

  PIN CON
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.0735 ;
  ANTENNAPARTIALMETALAREA 1.9443 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.6956 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10 0.69 10.34 1.03 ;
      RECT 8.95 0.79 10 1.02 ;
      RECT 9.1 2.91 9.58 3.25 ;
      RECT 8.95 1.82 9.1 3.25 ;
      RECT 8.72 0.79 8.95 3.48 ;
      RECT 8.18 1.27 8.72 1.61 ;
      RECT 8.32 3.25 8.72 3.48 ;
      RECT 8.12 3.25 8.32 4.155 ;
      RECT 8.09 3.25 8.12 4.21 ;
      RECT 7.78 3.87 8.09 4.21 ;
     END
  END CON

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.095 ;
  ANTENNAPARTIALMETALAREA 0.2501 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3409 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.23 2.405 14.305 2.635 ;
      RECT 14.02 2.105 14.23 2.635 ;
      RECT 14 1.995 14.02 2.635 ;
      RECT 13.68 1.995 14 2.335 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3608 ;
  ANTENNAPARTIALMETALAREA 0.242 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.113 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.93 1.75 7.23 2.1 ;
      RECT 6.615 1.75 6.93 2.185 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7452 ;
  ANTENNAPARTIALMETALAREA 0.231 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0282 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.875 2.11 1.295 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.58 -0.4 15.84 0.4 ;
      RECT 14.24 -0.4 14.58 1.655 ;
      RECT 14.16 -0.4 14.24 0.96 ;
      RECT 13.18 -0.4 14.16 0.4 ;
      RECT 12.84 -0.4 13.18 0.575 ;
      RECT 6.62 -0.4 12.84 0.4 ;
      RECT 6.28 -0.4 6.62 0.575 ;
      RECT 2.34 -0.4 6.28 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 1.225 -0.4 2 0.4 ;
      RECT 0.995 -0.4 1.225 0.67 ;
      RECT 0 -0.4 0.995 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.28 4.64 15.84 5.44 ;
      RECT 13.94 4.465 14.28 5.44 ;
      RECT 12.465 4.64 13.94 5.44 ;
      RECT 12.125 4.465 12.465 5.44 ;
      RECT 6.68 4.64 12.125 5.44 ;
      RECT 6.34 4.145 6.68 5.44 ;
      RECT 2.34 4.64 6.34 5.44 ;
      RECT 2 4.465 2.34 5.44 ;
      RECT 1.225 4.64 2 5.44 ;
      RECT 0.995 3.975 1.225 5.44 ;
      RECT 0 4.64 0.995 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.515 3.56 15.57 3.9 ;
      RECT 15.23 3.56 15.515 4.12 ;
      RECT 10.94 3.89 15.23 4.12 ;
      RECT 13.385 1.36 13.86 1.7 ;
      RECT 13.385 2.93 13.44 3.27 ;
      RECT 13.155 0.805 13.385 3.27 ;
      RECT 12.16 0.805 13.155 1.035 ;
      RECT 12.245 2.13 13.155 2.48 ;
      RECT 13.1 2.93 13.155 3.27 ;
      RECT 12.16 1.265 12.42 1.495 ;
      RECT 11.93 0.63 12.16 1.035 ;
      RECT 11.965 1.265 12.16 1.9 ;
      RECT 11.93 1.265 11.965 3.08 ;
      RECT 10.885 0.63 11.93 0.86 ;
      RECT 11.735 1.67 11.93 3.08 ;
      RECT 11.705 2.85 11.735 3.08 ;
      RECT 11.365 2.85 11.705 3.66 ;
      RECT 11.505 1.1 11.7 1.44 ;
      RECT 11.36 1.1 11.505 2.515 ;
      RECT 11.275 1.21 11.36 2.515 ;
      RECT 10.94 2.285 11.275 2.515 ;
      RECT 10.71 2.285 10.94 4.12 ;
      RECT 10.655 0.63 10.885 1.81 ;
      RECT 10.6 3.105 10.71 3.915 ;
      RECT 10.18 1.58 10.655 1.81 ;
      RECT 9.95 1.58 10.18 4.11 ;
      RECT 9.62 1.58 9.95 1.81 ;
      RECT 9.84 3.77 9.95 4.11 ;
      RECT 8.805 3.88 9.84 4.11 ;
      RECT 9.33 1.25 9.62 1.81 ;
      RECT 9.28 1.25 9.33 1.59 ;
      RECT 8.575 3.71 8.805 4.11 ;
      RECT 8.245 0.645 8.475 1.025 ;
      RECT 8.155 2.185 8.31 2.415 ;
      RECT 7.92 0.795 8.245 1.025 ;
      RECT 7.925 2.185 8.155 3.02 ;
      RECT 7.86 2.79 7.925 3.02 ;
      RECT 7.695 0.795 7.92 1.955 ;
      RECT 7.63 2.79 7.86 3.64 ;
      RECT 7.69 0.795 7.695 2.56 ;
      RECT 5.26 0.805 7.69 1.035 ;
      RECT 7.465 1.725 7.69 2.56 ;
      RECT 7.315 3.41 7.63 3.64 ;
      RECT 7.25 2.33 7.465 2.56 ;
      RECT 6.385 1.265 7.44 1.495 ;
      RECT 6.44 2.945 7.4 3.175 ;
      RECT 7.085 3.41 7.315 3.765 ;
      RECT 3.82 3.535 7.085 3.765 ;
      RECT 6.385 2.415 6.44 3.175 ;
      RECT 6.21 1.265 6.385 3.175 ;
      RECT 6.155 1.265 6.21 2.645 ;
      RECT 5.895 2.28 6.155 2.645 ;
      RECT 5.665 3.075 5.98 3.305 ;
      RECT 3.1 3.995 5.98 4.225 ;
      RECT 5.695 1.46 5.925 1.89 ;
      RECT 5.665 1.66 5.695 1.89 ;
      RECT 5.435 1.66 5.665 3.305 ;
      RECT 5.205 0.805 5.26 1.415 ;
      RECT 5.03 0.805 5.205 3.305 ;
      RECT 4.975 1.075 5.03 3.305 ;
      RECT 4.92 1.075 4.975 1.415 ;
      RECT 4.43 0.9 4.54 1.415 ;
      RECT 4.43 3.025 4.54 3.255 ;
      RECT 4.2 0.9 4.43 3.255 ;
      RECT 0.52 0.9 4.2 1.13 ;
      RECT 3.535 1.39 3.82 3.765 ;
      RECT 3.48 1.39 3.535 3.66 ;
      RECT 2.87 1.39 3.1 4.225 ;
      RECT 2.76 1.39 2.87 1.73 ;
      RECT 2.76 3.405 2.87 4.225 ;
      RECT 2.24 2.015 2.635 2.405 ;
      RECT 2.01 1.475 2.24 3.365 ;
      RECT 1.78 1.475 2.01 1.705 ;
      RECT 1.78 3.135 2.01 3.365 ;
      RECT 1.44 1.365 1.78 1.705 ;
      RECT 1.44 3.135 1.78 3.475 ;
      RECT 0.18 0.89 0.52 4.025 ;
  END
END AFHCONX4

MACRO AFHCONX2
  CLASS CORE ;
  FOREIGN AFHCONX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.52 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AFHCONX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2393 ;
  ANTENNAPARTIALMETALAREA 0.9832 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.4573 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.9 0.965 14.24 1.775 ;
      RECT 13.72 1.545 13.9 1.775 ;
      RECT 13.645 1.545 13.72 1.845 ;
      RECT 13.415 1.545 13.645 2.66 ;
      RECT 13.075 2.43 13.415 2.66 ;
      RECT 12.845 2.43 13.075 3.775 ;
     END
  END S

  PIN CON
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.888 ;
  ANTENNAPARTIALMETALAREA 1.0102 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.7753 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.95 1.845 9.025 2.075 ;
      RECT 8.72 1.325 8.95 3.195 ;
      RECT 8.68 1.325 8.72 1.61 ;
      RECT 8.59 2.965 8.72 3.195 ;
      RECT 8.34 1.27 8.68 1.61 ;
      RECT 8.36 2.965 8.59 3.535 ;
      RECT 8.265 3.305 8.36 3.535 ;
      RECT 8.035 3.305 8.265 4.15 ;
      RECT 7.78 3.92 8.035 4.15 ;
     END
  END CON

  PIN CI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5364 ;
  ANTENNAPARTIALMETALAREA 0.2226 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.007 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.04 1.82 12.46 2.35 ;
     END
  END CI

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3608 ;
  ANTENNAPARTIALMETALAREA 0.3249 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3091 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.74 1.805 7.12 2.66 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7434 ;
  ANTENNAPARTIALMETALAREA 0.2348 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0388 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.885 2.11 1.305 2.66 ;
      RECT 0.875 2.25 0.885 2.635 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 13.48 -0.4 14.52 0.4 ;
      RECT 13.14 -0.4 13.48 0.575 ;
      RECT 12.02 -0.4 13.14 0.4 ;
      RECT 11.68 -0.4 12.02 0.575 ;
      RECT 6.78 -0.4 11.68 0.4 ;
      RECT 6.44 -0.4 6.78 0.575 ;
      RECT 2.34 -0.4 6.44 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 1.28 -0.4 2 0.4 ;
      RECT 0.94 -0.4 1.28 0.635 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.37 4.64 14.52 5.44 ;
      RECT 12.03 4.465 12.37 5.44 ;
      RECT 11.145 4.64 12.03 5.44 ;
      RECT 10.805 4.465 11.145 5.44 ;
      RECT 6.68 4.64 10.805 5.44 ;
      RECT 6.34 4.145 6.68 5.44 ;
      RECT 2.34 4.64 6.34 5.44 ;
      RECT 2 4.465 2.34 5.44 ;
      RECT 1.28 4.64 2 5.44 ;
      RECT 0.94 4.185 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 13.515 2.9 13.745 4.235 ;
      RECT 9.87 4.005 13.515 4.235 ;
      RECT 12.44 0.765 12.78 1.575 ;
      RECT 11.725 1.055 12.44 1.285 ;
      RECT 11.725 1.8 11.75 3.775 ;
      RECT 11.52 0.805 11.725 3.775 ;
      RECT 11.495 0.805 11.52 2.085 ;
      RECT 11 0.805 11.495 1.035 ;
      RECT 11.39 1.725 11.495 2.085 ;
      RECT 11.15 1.265 11.26 1.495 ;
      RECT 10.92 1.265 11.15 1.78 ;
      RECT 10.77 0.63 11 1.035 ;
      RECT 10.645 1.55 10.92 1.78 ;
      RECT 9.725 0.63 10.77 0.86 ;
      RECT 10.415 1.55 10.645 3.66 ;
      RECT 10.185 1.09 10.54 1.32 ;
      RECT 10.33 3.43 10.415 3.66 ;
      RECT 10.1 3.43 10.33 3.775 ;
      RECT 9.955 1.09 10.185 3.2 ;
      RECT 9.87 2.97 9.955 3.2 ;
      RECT 9.64 2.97 9.87 4.235 ;
      RECT 9.495 0.63 9.725 2.735 ;
      RECT 9.28 3.885 9.64 4.115 ;
      RECT 9.41 2.505 9.495 2.735 ;
      RECT 9.18 2.505 9.41 3.655 ;
      RECT 9.05 3.425 9.18 3.655 ;
      RECT 8.86 3.425 9.05 3.995 ;
      RECT 8.82 3.425 8.86 4.105 ;
      RECT 8.52 3.765 8.82 4.105 ;
      RECT 8.35 0.645 8.69 1.035 ;
      RECT 8.13 2.185 8.44 2.415 ;
      RECT 8.08 0.805 8.35 1.035 ;
      RECT 7.9 2.185 8.13 3.075 ;
      RECT 7.85 0.805 8.08 1.955 ;
      RECT 7.805 2.845 7.9 3.075 ;
      RECT 5.42 0.805 7.85 1.035 ;
      RECT 7.67 1.725 7.85 1.955 ;
      RECT 7.575 2.845 7.805 3.69 ;
      RECT 7.44 1.725 7.67 2.615 ;
      RECT 6.51 1.265 7.6 1.495 ;
      RECT 6.795 3.46 7.575 3.69 ;
      RECT 7.115 2.89 7.345 3.23 ;
      RECT 6.51 2.89 7.115 3.12 ;
      RECT 6.565 3.46 6.795 3.765 ;
      RECT 3.82 3.535 6.565 3.765 ;
      RECT 6.28 1.265 6.51 3.12 ;
      RECT 5.95 2.335 6.28 2.565 ;
      RECT 5.72 2.92 5.98 3.15 ;
      RECT 3.1 3.995 5.98 4.225 ;
      RECT 5.72 1.46 5.925 1.89 ;
      RECT 5.695 1.46 5.72 3.15 ;
      RECT 5.49 1.66 5.695 3.15 ;
      RECT 5.26 0.805 5.42 1.36 ;
      RECT 5.19 0.805 5.26 1.415 ;
      RECT 5.15 3.075 5.26 3.305 ;
      RECT 5.15 1.075 5.19 1.415 ;
      RECT 4.92 1.075 5.15 3.305 ;
      RECT 4.425 0.865 4.54 1.415 ;
      RECT 4.425 3.075 4.54 3.305 ;
      RECT 4.195 0.865 4.425 3.305 ;
      RECT 0.52 0.865 4.195 1.095 ;
      RECT 3.535 1.39 3.82 3.765 ;
      RECT 3.48 1.39 3.535 3.66 ;
      RECT 2.87 1.39 3.1 4.225 ;
      RECT 2.76 1.39 2.87 1.73 ;
      RECT 2.76 3.405 2.87 4.225 ;
      RECT 2.24 2.015 2.635 2.405 ;
      RECT 2.01 1.475 2.24 3.26 ;
      RECT 1.78 1.475 2.01 1.705 ;
      RECT 1.78 3.03 2.01 3.26 ;
      RECT 1.44 1.365 1.78 1.705 ;
      RECT 1.44 3.03 1.78 3.37 ;
      RECT 0.465 0.765 0.52 1.575 ;
      RECT 0.235 0.765 0.465 4.02 ;
      RECT 0.18 0.765 0.235 1.575 ;
  END
END AFHCONX2

MACRO AFHCINX4
  CLASS CORE ;
  FOREIGN AFHCINX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.16 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.2658 ;
  ANTENNAPARTIALMETALAREA 0.9783 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7365 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.79 1.345 17.02 4.34 ;
      RECT 16.64 1.345 16.79 1.685 ;
      RECT 16.64 2.75 16.79 4.34 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 2.7685 ;
  ANTENNAPARTIALMETALAREA 1.8301 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.6532 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 11.65 1.29 11.88 1.685 ;
      RECT 10.775 1.29 11.65 1.52 ;
      RECT 10.925 2.865 11.155 3.24 ;
      RECT 10.895 3.01 10.925 3.24 ;
      RECT 10.665 3.01 10.895 3.775 ;
      RECT 10.495 1.29 10.775 1.54 ;
      RECT 9.77 3.545 10.665 3.775 ;
      RECT 10.225 1.29 10.495 1.63 ;
      RECT 9.995 1.29 10.225 2.305 ;
      RECT 9.77 2.075 9.995 2.305 ;
      RECT 9.76 2.075 9.77 3.775 ;
      RECT 9.54 2.075 9.76 3.78 ;
      RECT 9.38 2.38 9.54 3.78 ;
     END
  END CO

  PIN CIN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.0968 ;
  ANTENNAPARTIALMETALAREA 0.2373 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1077 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.68 2.38 15.7 2.66 ;
      RECT 15.34 1.995 15.68 2.66 ;
      RECT 15.32 2.38 15.34 2.66 ;
     END
  END CIN

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4716 ;
  ANTENNAPARTIALMETALAREA 0.2704 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1024 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.4 2.2 7.915 2.725 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7434 ;
  ANTENNAPARTIALMETALAREA 0.2327 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.36 2.17 1.835 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.345 -0.4 17.16 0.4 ;
      RECT 16.005 -0.4 16.345 0.965 ;
      RECT 15.025 -0.4 16.005 0.4 ;
      RECT 14.685 -0.4 15.025 0.575 ;
      RECT 7.945 -0.4 14.685 0.4 ;
      RECT 7.605 -0.4 7.945 0.575 ;
      RECT 2.34 -0.4 7.605 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 0.52 -0.4 2 0.4 ;
      RECT 0.18 -0.4 0.52 1.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 16.34 4.64 17.16 5.44 ;
      RECT 16 4.09 16.34 5.44 ;
      RECT 14.99 4.64 16 5.44 ;
      RECT 14.65 4.465 14.99 5.44 ;
      RECT 8.045 4.64 14.65 5.44 ;
      RECT 7.705 4.465 8.045 5.44 ;
      RECT 2.34 4.64 7.705 5.44 ;
      RECT 2 4.465 2.34 5.44 ;
      RECT 0.52 4.64 2 5.44 ;
      RECT 0.18 2.95 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 16.32 2.03 16.545 2.385 ;
      RECT 16.09 2.03 16.32 3.79 ;
      RECT 15.665 3.56 16.09 3.79 ;
      RECT 14.935 1.36 15.675 1.59 ;
      RECT 14.935 2.91 15.675 3.25 ;
      RECT 15.435 3.56 15.665 4.07 ;
      RECT 12.175 3.84 15.435 4.07 ;
      RECT 14.705 0.805 14.935 3.61 ;
      RECT 14.29 0.805 14.705 1.035 ;
      RECT 14.7 1.36 14.705 3.14 ;
      RECT 12.405 3.38 14.705 3.61 ;
      RECT 14.48 2.205 14.7 2.56 ;
      RECT 14.06 0.665 14.29 1.035 ;
      RECT 14.02 1.27 14.25 3.15 ;
      RECT 12.34 0.665 14.06 0.895 ;
      RECT 13.98 1.27 14.02 1.63 ;
      RECT 13.89 2.92 14.02 3.15 ;
      RECT 13.73 1.915 13.79 2.255 ;
      RECT 13.5 1.125 13.73 2.255 ;
      RECT 12.8 1.125 13.5 1.355 ;
      RECT 13.03 1.585 13.26 3.07 ;
      RECT 12.13 2.84 13.03 3.07 ;
      RECT 12.57 1.125 12.8 2.605 ;
      RECT 11.67 2.375 12.57 2.605 ;
      RECT 12.11 0.665 12.34 2.145 ;
      RECT 12.13 3.84 12.175 4.235 ;
      RECT 11.9 2.84 12.13 4.235 ;
      RECT 10.875 0.665 12.11 0.895 ;
      RECT 10.69 1.915 12.11 2.145 ;
      RECT 11.64 4.005 11.9 4.235 ;
      RECT 11.44 2.375 11.67 3.745 ;
      RECT 11.365 3.515 11.44 3.745 ;
      RECT 11.135 3.515 11.365 4.26 ;
      RECT 8.97 4.03 11.135 4.26 ;
      RECT 10.46 1.915 10.69 2.78 ;
      RECT 10.435 2.55 10.46 2.78 ;
      RECT 10.205 2.55 10.435 3.205 ;
      RECT 9.05 1.445 9.72 1.82 ;
      RECT 6.675 0.805 9.24 1.035 ;
      RECT 8.82 1.445 9.05 3.76 ;
      RECT 8.74 4.005 8.97 4.26 ;
      RECT 8.365 1.725 8.82 1.955 ;
      RECT 8.71 2.95 8.82 3.76 ;
      RECT 3.52 4.005 8.74 4.235 ;
      RECT 6.575 3.53 8.71 3.76 ;
      RECT 8.18 2.29 8.41 3.235 ;
      RECT 7.13 3.005 8.18 3.235 ;
      RECT 7.13 1.725 7.185 1.955 ;
      RECT 6.9 1.725 7.13 3.235 ;
      RECT 6.845 1.725 6.9 2.595 ;
      RECT 6.845 3.005 6.9 3.235 ;
      RECT 6.71 2.23 6.845 2.595 ;
      RECT 6.445 0.63 6.675 1.035 ;
      RECT 6.47 1.315 6.575 1.875 ;
      RECT 6.47 3.045 6.575 3.76 ;
      RECT 6.345 1.315 6.47 3.76 ;
      RECT 5.285 0.63 6.445 0.86 ;
      RECT 6.24 1.645 6.345 3.275 ;
      RECT 5.775 1.09 6.005 3.77 ;
      RECT 3.1 3.54 5.775 3.77 ;
      RECT 5.055 0.63 5.285 3.31 ;
      RECT 4.28 0.865 4.62 3.31 ;
      RECT 1.24 0.865 4.28 1.095 ;
      RECT 3.52 1.39 3.86 3.31 ;
      RECT 2.87 1.39 3.1 4.225 ;
      RECT 2.76 1.39 2.87 1.73 ;
      RECT 2.76 3.405 2.87 4.225 ;
      RECT 2.3 2.015 2.635 2.405 ;
      RECT 2.07 1.475 2.3 3.12 ;
      RECT 1.78 1.475 2.07 1.705 ;
      RECT 1.78 2.89 2.07 3.12 ;
      RECT 1.44 1.365 1.78 1.705 ;
      RECT 1.44 2.89 1.78 3.23 ;
      RECT 1.13 0.665 1.24 1.095 ;
      RECT 1.13 3.645 1.24 3.875 ;
      RECT 0.9 0.665 1.13 3.875 ;
  END
END AFHCINX4

MACRO AFHCINX2
  CLASS CORE ;
  FOREIGN AFHCINX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.84 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ AFHCINX4 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1412 ;
  ANTENNAPARTIALMETALAREA 0.9798 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.7365 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.47 1.345 15.7 4.34 ;
      RECT 15.32 1.345 15.47 1.685 ;
      RECT 15.32 2.74 15.47 4.34 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4653 ;
  ANTENNAPARTIALMETALAREA 0.9612 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.1499 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.225 1.11 10.495 1.45 ;
      RECT 9.995 1.11 10.225 2.455 ;
      RECT 9.77 2.225 9.995 2.455 ;
      RECT 9.54 2.225 9.77 3.91 ;
      RECT 9.43 2.94 9.54 3.91 ;
      RECT 9.38 2.94 9.43 3.22 ;
     END
  END CO

  PIN CIN
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5334 ;
  ANTENNAPARTIALMETALAREA 0.238 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1501 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.255 2.17 14.595 2.66 ;
      RECT 14 2.38 14.255 2.66 ;
     END
  END CIN

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.495 ;
  ANTENNAPARTIALMETALAREA 0.2151 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1925 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.595 1.82 7.78 2.1 ;
      RECT 7.365 1.82 7.595 2.53 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7434 ;
  ANTENNAPARTIALMETALAREA 0.2327 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0229 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.36 2.17 1.835 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 15.025 -0.4 15.84 0.4 ;
      RECT 14.685 -0.4 15.025 1.055 ;
      RECT 13.705 -0.4 14.685 0.4 ;
      RECT 13.365 -0.4 13.705 0.575 ;
      RECT 7.93 -0.4 13.365 0.4 ;
      RECT 7.59 -0.4 7.93 0.575 ;
      RECT 2.34 -0.4 7.59 0.4 ;
      RECT 2 -0.4 2.34 0.575 ;
      RECT 0.52 -0.4 2 0.4 ;
      RECT 0.18 -0.4 0.52 1.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 14.9 4.64 15.84 5.44 ;
      RECT 14.56 3.995 14.9 5.44 ;
      RECT 12.895 4.64 14.56 5.44 ;
      RECT 12.555 4.465 12.895 5.44 ;
      RECT 8.205 4.64 12.555 5.44 ;
      RECT 7.865 4.465 8.205 5.44 ;
      RECT 2.34 4.64 7.865 5.44 ;
      RECT 2 4.465 2.34 5.44 ;
      RECT 0.52 4.64 2 5.44 ;
      RECT 0.18 2.95 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 15.055 2.03 15.225 2.385 ;
      RECT 14.825 2.03 15.055 3.73 ;
      RECT 13.355 3.5 14.825 3.73 ;
      RECT 13.73 1.36 14.355 1.7 ;
      RECT 13.84 2.91 14.18 3.25 ;
      RECT 13.73 2.91 13.84 3.14 ;
      RECT 13.5 0.805 13.73 3.14 ;
      RECT 13.005 0.805 13.5 1.035 ;
      RECT 13.125 2.555 13.5 2.895 ;
      RECT 13.125 3.5 13.355 4.105 ;
      RECT 11.615 3.875 13.125 4.105 ;
      RECT 12.775 0.665 13.005 1.035 ;
      RECT 12.66 1.27 12.89 3.525 ;
      RECT 10.96 0.665 12.775 0.895 ;
      RECT 12.08 3.295 12.66 3.525 ;
      RECT 12.185 1.125 12.415 2.455 ;
      RECT 11.42 1.125 12.185 1.355 ;
      RECT 11.85 3.295 12.08 3.64 ;
      RECT 11.71 1.585 11.94 2.97 ;
      RECT 11.615 2.74 11.71 2.97 ;
      RECT 11.385 2.74 11.615 4.105 ;
      RECT 11.19 1.125 11.42 2.49 ;
      RECT 11.125 3.695 11.385 4.105 ;
      RECT 11.145 2.26 11.19 2.49 ;
      RECT 10.915 2.26 11.145 3.415 ;
      RECT 10.73 0.665 10.96 1.985 ;
      RECT 10.895 3.185 10.915 3.415 ;
      RECT 10.665 3.185 10.895 4.385 ;
      RECT 10.685 1.755 10.73 1.985 ;
      RECT 10.455 1.755 10.685 2.925 ;
      RECT 9.13 4.155 10.665 4.385 ;
      RECT 10.435 2.695 10.455 2.925 ;
      RECT 10.205 2.695 10.435 3.91 ;
      RECT 9.49 1.23 9.72 1.835 ;
      RECT 8.995 1.605 9.49 1.835 ;
      RECT 5.34 0.805 9.23 1.035 ;
      RECT 8.9 4.005 9.13 4.385 ;
      RECT 8.995 2.965 9.05 3.775 ;
      RECT 8.765 1.605 8.995 3.775 ;
      RECT 4.775 4.005 8.9 4.235 ;
      RECT 8.35 1.605 8.765 1.835 ;
      RECT 8.71 2.965 8.765 3.775 ;
      RECT 6.465 3.455 8.71 3.685 ;
      RECT 8.205 2.275 8.435 3.16 ;
      RECT 7.115 2.93 8.205 3.16 ;
      RECT 6.885 1.545 7.115 3.16 ;
      RECT 6.695 2.15 6.885 2.55 ;
      RECT 6.465 1.355 6.535 1.725 ;
      RECT 6.235 1.355 6.465 3.685 ;
      RECT 5.775 1.29 6.005 3.77 ;
      RECT 3.1 3.485 5.775 3.715 ;
      RECT 5 0.805 5.34 3.245 ;
      RECT 4.545 3.945 4.775 4.235 ;
      RECT 4.28 0.865 4.62 3.245 ;
      RECT 3.52 3.945 4.545 4.175 ;
      RECT 1.24 0.865 4.28 1.095 ;
      RECT 3.52 1.39 3.86 3.245 ;
      RECT 2.87 1.39 3.1 4.225 ;
      RECT 2.76 1.39 2.87 1.73 ;
      RECT 2.76 3.405 2.87 4.225 ;
      RECT 2.3 2.015 2.635 2.405 ;
      RECT 2.07 1.475 2.3 3.12 ;
      RECT 1.78 1.475 2.07 1.705 ;
      RECT 1.78 2.89 2.07 3.12 ;
      RECT 1.44 1.365 1.78 1.705 ;
      RECT 1.44 2.89 1.78 3.23 ;
      RECT 1.13 0.665 1.24 1.095 ;
      RECT 1.13 3.645 1.24 3.875 ;
      RECT 0.9 0.665 1.13 3.875 ;
  END
END AFHCINX2

MACRO CMPR42X2
  CLASS CORE ;
  FOREIGN CMPR42X2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 26.4 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.3968 ;
  ANTENNAPARTIALMETALAREA 0.86 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4344 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 26.185 0.765 26.22 1.575 ;
      RECT 26.185 2.38 26.22 3.555 ;
      RECT 25.955 0.765 26.185 3.555 ;
      RECT 25.88 0.765 25.955 1.575 ;
      RECT 25.88 2.38 25.955 3.555 ;
     END
  END S

  PIN ICO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.4256 ;
  ANTENNAPARTIALMETALAREA 0.7888 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.2648 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.4 0.945 0.52 1.755 ;
      RECT 0.4 2.745 0.52 3.555 ;
      RECT 0.18 0.945 0.4 3.555 ;
      RECT 0.17 1.235 0.18 3.265 ;
     END
  END ICO

  PIN ICI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4662 ;
  ANTENNAPARTIALMETALAREA 0.2254 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.895 1.875 23.045 2.105 ;
      RECT 22.665 1.285 22.895 2.105 ;
      RECT 22.655 1.285 22.665 1.515 ;
     END
  END ICI

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9828 ;
  ANTENNAPARTIALMETALAREA 0.7911 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.8902 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.945 1.985 17.47 2.215 ;
      RECT 16.715 1.845 16.945 2.24 ;
      RECT 15.06 2.01 16.715 2.24 ;
      RECT 14.83 2.01 15.06 2.665 ;
      RECT 14.62 2.435 14.83 2.665 ;
     END
  END D

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.1896 ;
  ANTENNAPARTIALMETALAREA 0.7211 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4874 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.73 2.965 20.905 3.195 ;
      RECT 20.52 1.265 20.73 3.36 ;
      RECT 20.5 1.265 20.52 3.445 ;
      RECT 20.115 1.265 20.5 1.495 ;
      RECT 20.18 3.105 20.5 3.445 ;
     END
  END CO

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.9054 ;
  ANTENNAPARTIALMETALAREA 3.4701 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 16.0802 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.195 4.175 17.25 4.405 ;
      RECT 16.285 4.175 17.195 4.41 ;
      RECT 16.055 4.085 16.285 4.41 ;
      RECT 14.405 4.085 16.055 4.315 ;
      RECT 14.175 4.005 14.405 4.315 ;
      RECT 13.375 4.005 14.175 4.235 ;
      RECT 13.145 4.005 13.375 4.41 ;
      RECT 10.425 4.18 13.145 4.41 ;
      RECT 10.195 4.005 10.425 4.41 ;
      RECT 9.39 4.005 10.195 4.235 ;
      RECT 9.16 4.005 9.39 4.405 ;
      RECT 7.06 4.175 9.16 4.405 ;
      RECT 6.83 4.005 7.06 4.405 ;
      RECT 4.175 4.005 6.83 4.235 ;
      RECT 3.895 4.005 4.175 4.34 ;
      RECT 3.665 4.005 3.895 4.41 ;
      RECT 3.35 4.18 3.665 4.41 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.4742 ;
  ANTENNAPARTIALMETALAREA 1.9932 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.3333 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.01 2.525 8.45 2.755 ;
      RECT 7.78 2.525 8.01 2.985 ;
      RECT 6.565 2.755 7.78 2.985 ;
      RECT 6.335 2.755 6.565 3.625 ;
      RECT 5.295 3.395 6.335 3.625 ;
      RECT 5.295 2.265 5.35 2.495 ;
      RECT 5.065 2.265 5.295 3.625 ;
      RECT 3.82 2.265 5.065 2.495 ;
      RECT 3.44 2.265 3.82 2.635 ;
      RECT 2.07 2.265 3.44 2.495 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.3248 ;
  ANTENNAPARTIALMETALAREA 1.3006 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 6.2381 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.765 1.8 6.515 2.03 ;
      RECT 1.69 1.8 1.765 2.075 ;
      RECT 1.535 1.8 1.69 2.415 ;
      RECT 1.46 1.845 1.535 2.415 ;
      RECT 1.245 2.185 1.46 2.415 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 25.46 -0.4 26.4 0.4 ;
      RECT 25.12 -0.4 25.46 0.575 ;
      RECT 22.655 -0.4 25.12 0.4 ;
      RECT 22.315 -0.4 22.655 0.575 ;
      RECT 21.45 -0.4 22.315 0.4 ;
      RECT 21.11 -0.4 21.45 0.575 ;
      RECT 17.315 -0.4 21.11 0.4 ;
      RECT 16.975 -0.4 17.315 0.575 ;
      RECT 13.205 -0.4 16.975 0.4 ;
      RECT 12.865 -0.4 13.205 0.575 ;
      RECT 9.65 -0.4 12.865 0.4 ;
      RECT 9.31 -0.4 9.65 0.575 ;
      RECT 6.85 -0.4 9.31 0.4 ;
      RECT 6.51 -0.4 6.85 0.575 ;
      RECT 5.38 -0.4 6.51 0.4 ;
      RECT 5.04 -0.4 5.38 0.575 ;
      RECT 3.86 -0.4 5.04 0.4 ;
      RECT 3.52 -0.4 3.86 0.575 ;
      RECT 1.28 -0.4 3.52 0.4 ;
      RECT 0.94 -0.4 1.28 0.575 ;
      RECT 0 -0.4 0.94 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 25.46 4.64 26.4 5.44 ;
      RECT 25.405 4.465 25.46 5.44 ;
      RECT 25.175 3.32 25.405 5.44 ;
      RECT 25.12 4.465 25.175 5.44 ;
      RECT 22.405 4.64 25.12 5.44 ;
      RECT 22.065 4.465 22.405 5.44 ;
      RECT 17.71 4.64 22.065 5.44 ;
      RECT 17.48 3.71 17.71 5.44 ;
      RECT 17.25 3.71 17.48 3.94 ;
      RECT 13.945 4.64 17.48 5.44 ;
      RECT 16.91 3.13 17.25 3.94 ;
      RECT 13.605 4.465 13.945 5.44 ;
      RECT 9.96 4.64 13.605 5.44 ;
      RECT 9.62 4.465 9.96 5.44 ;
      RECT 6.6 4.64 9.62 5.44 ;
      RECT 6.26 4.465 6.6 5.44 ;
      RECT 5.54 4.64 6.26 5.44 ;
      RECT 5.2 4.465 5.54 5.44 ;
      RECT 1.28 4.64 5.2 5.44 ;
      RECT 0.94 3.84 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 25.43 1.92 25.725 2.15 ;
      RECT 25.2 0.805 25.43 3.09 ;
      RECT 23.795 0.805 25.2 1.035 ;
      RECT 24.945 2.86 25.2 3.09 ;
      RECT 24.74 1.265 24.97 2.63 ;
      RECT 24.89 2.86 24.945 4.19 ;
      RECT 24.715 2.86 24.89 4.25 ;
      RECT 23.55 1.265 24.74 1.495 ;
      RECT 24.485 2.4 24.74 2.63 ;
      RECT 24.66 3.96 24.715 4.25 ;
      RECT 23.885 4.02 24.66 4.25 ;
      RECT 23.505 1.725 24.51 1.955 ;
      RECT 24.43 2.4 24.485 3.405 ;
      RECT 24.255 2.4 24.43 3.79 ;
      RECT 24.2 3.175 24.255 3.79 ;
      RECT 23.165 3.56 24.2 3.79 ;
      RECT 23.97 2.58 24.025 2.945 ;
      RECT 23.795 2.58 23.97 3.33 ;
      RECT 23.545 4.02 23.885 4.36 ;
      RECT 23.74 2.715 23.795 3.33 ;
      RECT 21.835 3.1 23.74 3.33 ;
      RECT 23.32 0.8 23.55 1.495 ;
      RECT 23.275 1.725 23.505 2.775 ;
      RECT 23.075 0.8 23.32 1.03 ;
      RECT 22.35 2.545 23.275 2.775 ;
      RECT 23.055 3.56 23.165 3.92 ;
      RECT 22.88 3.56 23.055 4.235 ;
      RECT 22.825 3.58 22.88 4.235 ;
      RECT 21.65 4.005 22.825 4.235 ;
      RECT 22.12 0.805 22.35 2.775 ;
      RECT 21.25 0.805 22.12 1.035 ;
      RECT 21.82 1.43 21.835 3.33 ;
      RECT 21.73 1.375 21.82 3.33 ;
      RECT 21.605 1.375 21.73 3.685 ;
      RECT 21.42 4.005 21.65 4.41 ;
      RECT 21.48 1.375 21.605 1.715 ;
      RECT 21.5 2.795 21.605 3.685 ;
      RECT 21.19 3.455 21.5 3.685 ;
      RECT 19.58 4.18 21.42 4.41 ;
      RECT 21.25 1.945 21.375 2.37 ;
      RECT 21.145 0.805 21.25 2.37 ;
      RECT 20.96 3.455 21.19 3.95 ;
      RECT 21.02 0.805 21.145 2.175 ;
      RECT 20.37 0.805 21.02 1.035 ;
      RECT 19.81 3.72 20.96 3.95 ;
      RECT 20.14 0.63 20.37 1.035 ;
      RECT 20.04 1.725 20.27 2.875 ;
      RECT 18.48 0.63 20.14 0.86 ;
      RECT 19.715 1.725 20.04 1.955 ;
      RECT 19.78 2.645 20.04 2.875 ;
      RECT 19.115 2.185 19.81 2.415 ;
      RECT 19.58 2.645 19.78 3.475 ;
      RECT 19.485 1.13 19.715 1.955 ;
      RECT 19.55 2.645 19.58 4.41 ;
      RECT 19.44 3.135 19.55 4.41 ;
      RECT 19.375 1.13 19.485 1.47 ;
      RECT 19.35 3.245 19.44 4.41 ;
      RECT 19.06 2 19.115 3.395 ;
      RECT 18.94 2 19.06 3.975 ;
      RECT 18.885 1.105 18.94 3.975 ;
      RECT 18.71 1.105 18.885 2.23 ;
      RECT 18.72 3.165 18.885 3.975 ;
      RECT 18.48 2.505 18.655 2.92 ;
      RECT 18.425 0.63 18.48 2.92 ;
      RECT 18.25 0.63 18.425 2.735 ;
      RECT 18 3.16 18.34 3.97 ;
      RECT 18.18 0.63 18.25 1.035 ;
      RECT 16.58 0.805 18.18 1.035 ;
      RECT 17.95 1.265 18.02 1.985 ;
      RECT 17.95 3.16 18 3.39 ;
      RECT 17.79 1.265 17.95 3.39 ;
      RECT 17.72 1.755 17.79 3.39 ;
      RECT 17.65 2.47 17.72 3.39 ;
      RECT 15.29 2.47 17.65 2.7 ;
      RECT 16.35 0.63 16.58 1.035 ;
      RECT 16.29 1.27 16.555 1.5 ;
      RECT 13.68 0.63 16.35 0.86 ;
      RECT 16.06 1.27 16.29 1.78 ;
      RECT 14.225 3.085 16.16 3.315 ;
      RECT 14.6 1.55 16.06 1.78 ;
      RECT 14.14 1.09 15.735 1.32 ;
      RECT 13.7 3.545 15.44 3.775 ;
      RECT 14.37 1.55 14.6 1.955 ;
      RECT 14.325 1.725 14.37 1.955 ;
      RECT 14.225 1.725 14.325 2.4 ;
      RECT 14.095 1.725 14.225 3.315 ;
      RECT 13.91 1.09 14.14 1.495 ;
      RECT 13.995 2.115 14.095 3.315 ;
      RECT 13.885 2.115 13.995 2.455 ;
      RECT 12.455 1.265 13.91 1.495 ;
      RECT 13.47 3.005 13.7 3.775 ;
      RECT 13.45 0.63 13.68 1.035 ;
      RECT 12.71 3.005 13.47 3.235 ;
      RECT 11.985 0.805 13.45 1.035 ;
      RECT 12.915 3.465 13.24 3.695 ;
      RECT 12.685 3.465 12.915 3.95 ;
      RECT 12.455 2.89 12.71 3.235 ;
      RECT 10.885 3.72 12.685 3.95 ;
      RECT 12.225 1.265 12.455 3.49 ;
      RECT 12.215 1.265 12.225 1.625 ;
      RECT 11.35 3.26 12.225 3.49 ;
      RECT 11.985 1.98 11.995 3.03 ;
      RECT 11.765 0.805 11.985 3.03 ;
      RECT 11.755 0.805 11.765 2.21 ;
      RECT 11.645 2.8 11.765 3.03 ;
      RECT 11.315 1.21 11.755 1.495 ;
      RECT 11.295 1.745 11.525 2.12 ;
      RECT 11.12 2.56 11.35 3.49 ;
      RECT 10.975 1.155 11.315 1.495 ;
      RECT 10.46 1.745 11.295 1.975 ;
      RECT 10.855 2.56 11.12 2.79 ;
      RECT 10.655 3.545 10.885 3.95 ;
      RECT 10.625 2.21 10.855 2.79 ;
      RECT 10.34 3.02 10.725 3.25 ;
      RECT 9.745 3.545 10.655 3.775 ;
      RECT 10.34 1.155 10.46 1.975 ;
      RECT 10.12 1.155 10.34 3.25 ;
      RECT 10.11 1.21 10.12 3.25 ;
      RECT 9.515 0.935 9.745 3.775 ;
      RECT 8.33 0.935 9.515 1.165 ;
      RECT 8.93 3.545 9.515 3.775 ;
      RECT 8.93 1.395 9.16 2.765 ;
      RECT 7.61 1.395 8.93 1.625 ;
      RECT 8.91 2.535 8.93 2.765 ;
      RECT 8.7 3.545 8.93 3.945 ;
      RECT 8.68 2.535 8.91 3.24 ;
      RECT 7.55 1.855 8.7 2.085 ;
      RECT 7.74 3.715 8.7 3.945 ;
      RECT 8.47 3.01 8.68 3.24 ;
      RECT 8.24 3.01 8.47 3.485 ;
      RECT 7.99 0.825 8.33 1.165 ;
      RECT 7.02 3.255 8.24 3.485 ;
      RECT 7.38 1.02 7.61 1.625 ;
      RECT 7.32 1.855 7.55 2.525 ;
      RECT 7.27 1.02 7.38 1.36 ;
      RECT 6.975 2.295 7.32 2.525 ;
      RECT 6.745 1.34 6.975 2.525 ;
      RECT 5.98 1.34 6.745 1.57 ;
      RECT 6.1 2.295 6.745 2.525 ;
      RECT 5.87 2.295 6.1 3.155 ;
      RECT 5.745 1.12 5.98 1.57 ;
      RECT 5.76 2.815 5.87 3.155 ;
      RECT 5.64 1.12 5.745 1.46 ;
      RECT 4.44 2.875 4.78 3.685 ;
      RECT 4.565 0.865 4.62 1.205 ;
      RECT 4.28 0.865 4.565 1.32 ;
      RECT 3.32 3.38 4.44 3.61 ;
      RECT 3.32 1.09 4.28 1.32 ;
      RECT 3.035 1.09 3.32 1.57 ;
      RECT 2.98 3.325 3.32 3.665 ;
      RECT 2.98 1.23 3.035 1.57 ;
      RECT 2.26 1.15 2.6 1.49 ;
      RECT 2.26 3.325 2.6 3.665 ;
      RECT 0.98 1.205 2.26 1.435 ;
      RECT 0.98 3.38 2.26 3.61 ;
      RECT 0.75 1.205 0.98 3.61 ;
      RECT 0.63 2.175 0.75 2.515 ;
  END
END CMPR42X2

MACRO CMPR42X1
  CLASS CORE ;
  FOREIGN CMPR42X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 22.44 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ CMPR42X2 ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7485 ;
  ANTENNAPARTIALMETALAREA 0.7647 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.1535 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 22.22 1.175 22.265 3.265 ;
      RECT 22.035 1.12 22.22 3.555 ;
      RECT 21.88 1.12 22.035 1.46 ;
      RECT 21.92 2.38 22.035 3.555 ;
      RECT 21.88 2.745 21.92 3.555 ;
     END
  END S

  PIN ICO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.744 ;
  ANTENNAPARTIALMETALAREA 0.6405 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8302 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.4 1.355 0.52 1.695 ;
      RECT 0.4 2.745 0.52 3.555 ;
      RECT 0.18 1.355 0.4 3.555 ;
      RECT 0.17 1.41 0.18 3.265 ;
     END
  END ICO

  PIN ICI
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.1728 ;
  ANTENNAPARTIALMETALAREA 0.2666 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2826 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 19.055 2.375 19.585 2.66 ;
      RECT 18.715 2.32 19.055 2.66 ;
     END
  END ICI

  PIN D
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4428 ;
  ANTENNAPARTIALMETALAREA 0.4394 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.0511 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.34 1.8 14 2.14 ;
      RECT 12.845 1.8 13.34 2.03 ;
      RECT 12.615 1.59 12.845 2.03 ;
     END
  END D

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.7192 ;
  ANTENNAPARTIALMETALAREA 0.5209 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4115 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.94 1.37 16.995 1.845 ;
      RECT 16.945 2.635 16.995 3.08 ;
      RECT 16.94 2.635 16.945 3.195 ;
      RECT 16.715 1.37 16.94 3.195 ;
      RECT 16.71 1.37 16.715 3.08 ;
      RECT 16.655 1.37 16.71 1.845 ;
      RECT 16.655 2.635 16.71 3.08 ;
     END
  END CO

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4428 ;
  ANTENNAPARTIALMETALAREA 2.5663 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.6865 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.06 3.95 13.09 4.29 ;
      RECT 12.75 3.5 13.06 4.29 ;
      RECT 12.68 3.5 12.75 4.235 ;
      RECT 6.305 4.005 12.68 4.235 ;
      RECT 6.075 4.005 6.305 4.41 ;
      RECT 3.03 4.18 6.075 4.41 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7164 ;
  ANTENNAPARTIALMETALAREA 0.4427 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.2843 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.745 1.88 3.99 2.11 ;
      RECT 3.515 1.845 3.745 2.11 ;
      RECT 2.1 1.88 3.515 2.11 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.6048 ;
  ANTENNAPARTIALMETALAREA 1.0292 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.8124 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.65 1.985 4.76 2.325 ;
      RECT 4.42 1.985 4.65 2.57 ;
      RECT 1.765 2.34 4.42 2.57 ;
      RECT 1.535 1.845 1.765 2.57 ;
      RECT 1.3 2.1 1.535 2.44 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 21.42 -0.4 22.44 0.4 ;
      RECT 21.08 -0.4 21.42 0.575 ;
      RECT 18.225 -0.4 21.08 0.4 ;
      RECT 17.415 -0.4 18.225 0.575 ;
      RECT 13.85 -0.4 17.415 0.4 ;
      RECT 13.51 -0.4 13.85 0.575 ;
      RECT 10.66 -0.4 13.51 0.4 ;
      RECT 10.32 -0.4 10.66 0.575 ;
      RECT 7.78 -0.4 10.32 0.4 ;
      RECT 7.44 -0.4 7.78 0.575 ;
      RECT 5.02 -0.4 7.44 0.4 ;
      RECT 4.68 -0.4 5.02 1.275 ;
      RECT 2.72 -0.4 4.68 0.4 ;
      RECT 2.38 -0.4 2.72 0.575 ;
      RECT 1.12 -0.4 2.38 0.4 ;
      RECT 0.78 -0.4 1.12 0.575 ;
      RECT 0 -0.4 0.78 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 21.655 4.64 22.44 5.44 ;
      RECT 21.315 4.465 21.655 5.44 ;
      RECT 18.775 4.64 21.315 5.44 ;
      RECT 18.435 3.81 18.775 5.44 ;
      RECT 17.755 4.64 18.435 5.44 ;
      RECT 17.415 4.465 17.755 5.44 ;
      RECT 13.66 4.64 17.415 5.44 ;
      RECT 13.32 2.885 13.66 5.44 ;
      RECT 11.06 4.64 13.32 5.44 ;
      RECT 10.72 4.465 11.06 5.44 ;
      RECT 7.58 4.64 10.72 5.44 ;
      RECT 7.24 4.465 7.58 5.44 ;
      RECT 2.8 4.64 7.24 5.44 ;
      RECT 4.925 3.41 4.98 3.75 ;
      RECT 4.64 3.41 4.925 3.95 ;
      RECT 2.8 3.72 4.64 3.95 ;
      RECT 2.57 3.72 2.8 5.44 ;
      RECT 2.46 4.465 2.57 5.44 ;
      RECT 1.28 4.64 2.46 5.44 ;
      RECT 0.94 4.465 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 21.65 1.805 21.805 2.145 ;
      RECT 21.42 1.555 21.65 4.04 ;
      RECT 20.795 1.555 21.42 1.785 ;
      RECT 20.295 3.81 21.42 4.04 ;
      RECT 20.98 2.015 21.135 2.355 ;
      RECT 20.75 2.015 20.98 3.58 ;
      RECT 20.565 0.785 20.795 1.785 ;
      RECT 20.32 2.015 20.75 2.245 ;
      RECT 19.535 3.35 20.75 3.58 ;
      RECT 19.72 0.785 20.565 1.015 ;
      RECT 20.18 2.78 20.52 3.12 ;
      RECT 20.09 1.245 20.32 2.245 ;
      RECT 19.955 3.81 20.295 4.15 ;
      RECT 18.365 2.89 20.18 3.12 ;
      RECT 19.26 1.245 20.09 1.475 ;
      RECT 18.365 1.705 19.61 1.935 ;
      RECT 19.195 3.35 19.535 3.79 ;
      RECT 19.03 0.76 19.26 1.475 ;
      RECT 17.955 3.35 19.195 3.58 ;
      RECT 18.92 0.76 19.03 1.1 ;
      RECT 18.135 1.375 18.365 3.12 ;
      RECT 18.015 1.375 18.135 1.715 ;
      RECT 18.015 2.74 18.135 3.12 ;
      RECT 17.48 2.89 18.015 3.12 ;
      RECT 17.725 3.35 17.955 4.145 ;
      RECT 17.785 2.03 17.905 2.37 ;
      RECT 17.555 0.805 17.785 2.37 ;
      RECT 17.075 3.915 17.725 4.145 ;
      RECT 17.05 0.805 17.555 1.035 ;
      RECT 17.25 2.89 17.48 3.685 ;
      RECT 16.615 3.455 17.25 3.685 ;
      RECT 16.845 3.915 17.075 4.38 ;
      RECT 16.82 0.63 17.05 1.035 ;
      RECT 15.895 4.15 16.845 4.38 ;
      RECT 14.92 0.63 16.82 0.86 ;
      RECT 16.385 3.455 16.615 3.92 ;
      RECT 16.125 3.69 16.385 3.92 ;
      RECT 16.035 1.105 16.235 1.445 ;
      RECT 15.895 1.105 16.035 3.225 ;
      RECT 15.805 1.105 15.895 4.38 ;
      RECT 15.665 2.885 15.805 4.38 ;
      RECT 15.38 4.065 15.435 4.405 ;
      RECT 15.15 1.105 15.38 4.405 ;
      RECT 14.975 2.955 15.15 3.295 ;
      RECT 15.095 4.065 15.15 4.405 ;
      RECT 14.69 0.63 14.92 2.695 ;
      RECT 13.28 0.805 14.69 1.035 ;
      RECT 14.42 1.32 14.46 2.6 ;
      RECT 14.23 1.32 14.42 3.295 ;
      RECT 14.12 1.32 14.23 1.55 ;
      RECT 14.08 2.37 14.23 3.295 ;
      RECT 12.66 2.37 14.08 2.6 ;
      RECT 13.05 0.63 13.28 1.035 ;
      RECT 11.145 0.63 13.05 0.86 ;
      RECT 12.56 2.83 12.9 3.17 ;
      RECT 12.385 1.09 12.82 1.32 ;
      RECT 12.32 2.26 12.66 2.6 ;
      RECT 11.18 2.83 12.56 3.06 ;
      RECT 12.155 1.09 12.385 1.955 ;
      RECT 11.84 3.295 12.18 3.635 ;
      RECT 11.18 1.725 12.155 1.955 ;
      RECT 11.695 1.09 11.925 1.495 ;
      RECT 10.36 3.295 11.84 3.525 ;
      RECT 10.385 1.265 11.695 1.495 ;
      RECT 10.95 1.725 11.18 3.06 ;
      RECT 10.915 0.63 11.145 1.035 ;
      RECT 10.84 2.26 10.95 2.6 ;
      RECT 9.53 0.805 10.915 1.035 ;
      RECT 10.385 1.89 10.44 2.23 ;
      RECT 10.36 1.265 10.385 2.23 ;
      RECT 10.155 1.265 10.36 3.695 ;
      RECT 9.82 1.265 10.155 1.495 ;
      RECT 10.13 1.89 10.155 3.695 ;
      RECT 10.1 1.89 10.13 2.23 ;
      RECT 10.02 2.885 10.13 3.695 ;
      RECT 9.53 2.885 9.64 3.695 ;
      RECT 9.3 0.805 9.53 3.695 ;
      RECT 9.1 1.155 9.3 1.495 ;
      RECT 7.775 3.545 8.88 3.775 ;
      RECT 8.53 1.155 8.575 1.495 ;
      RECT 8.39 0.63 8.53 1.495 ;
      RECT 8.345 0.63 8.39 3.075 ;
      RECT 8.19 0.63 8.345 3.13 ;
      RECT 8.16 1.21 8.19 3.13 ;
      RECT 8.005 2.79 8.16 3.13 ;
      RECT 7.775 2.22 7.93 2.56 ;
      RECT 7.545 1.09 7.775 3.775 ;
      RECT 6.46 1.09 7.545 1.32 ;
      RECT 6.46 3.545 7.545 3.775 ;
      RECT 7.15 1.985 7.26 2.325 ;
      RECT 6.92 1.775 7.15 3.06 ;
      RECT 5.74 1.775 6.92 2.005 ;
      RECT 5.685 2.83 6.92 3.06 ;
      RECT 6.12 0.98 6.46 1.32 ;
      RECT 6.175 3.295 6.46 3.775 ;
      RECT 6.12 3.295 6.175 3.635 ;
      RECT 5.64 2.26 5.98 2.6 ;
      RECT 5.51 0.955 5.74 2.005 ;
      RECT 5.455 2.83 5.685 3.675 ;
      RECT 5.22 2.315 5.64 2.6 ;
      RECT 5.4 0.955 5.51 1.295 ;
      RECT 4.99 1.525 5.22 3.16 ;
      RECT 4.45 1.525 4.99 1.755 ;
      RECT 4.18 2.93 4.99 3.16 ;
      RECT 4.22 1.145 4.45 1.755 ;
      RECT 3.88 1.035 4.22 1.375 ;
      RECT 3.84 2.93 4.18 3.275 ;
      RECT 3.41 1.235 3.52 1.575 ;
      RECT 3.37 2.92 3.48 3.26 ;
      RECT 3.18 0.805 3.41 1.575 ;
      RECT 3.14 2.92 3.37 3.49 ;
      RECT 1.92 0.805 3.18 1.035 ;
      RECT 2.04 3.26 3.14 3.49 ;
      RECT 0.98 2.8 2.76 3.03 ;
      RECT 2.38 1.295 2.72 1.635 ;
      RECT 0.98 1.35 2.38 1.58 ;
      RECT 1.81 3.26 2.04 4.345 ;
      RECT 1.635 0.63 1.92 1.035 ;
      RECT 1.7 4.005 1.81 4.345 ;
      RECT 1.58 0.63 1.635 0.97 ;
      RECT 0.75 1.35 0.98 3.03 ;
      RECT 0.63 2.03 0.75 2.37 ;
  END
END CMPR42X1

MACRO CMPR32X1
  CLASS CORE ;
  FOREIGN CMPR32X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.86 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.7191 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.0157 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.57 1.285 13.645 1.515 ;
      RECT 13.46 1.285 13.57 1.845 ;
      RECT 13.46 2.635 13.57 3.605 ;
      RECT 13.23 1.285 13.46 3.605 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.732 ;
  ANTENNAPARTIALMETALAREA 0.5743 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.6235 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.005 2.38 12.325 2.66 ;
      RECT 11.985 1.43 12.005 2.66 ;
      RECT 11.755 1.43 11.985 3.135 ;
      RECT 11.665 1.43 11.755 1.77 ;
      RECT 11.645 2.795 11.755 3.135 ;
     END
  END CO

  PIN C
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3816 ;
  ANTENNAPARTIALMETALAREA 0.5213 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.4221 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.22 1.82 9.485 2.05 ;
      RECT 8.99 1.82 9.22 3.22 ;
      RECT 8.6 2.865 8.99 3.22 ;
     END
  END C

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5424 ;
  ANTENNAPARTIALMETALAREA 0.2214 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.2084 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.445 2.04 0.76 2.38 ;
      RECT 0.42 2.04 0.445 2.635 ;
      RECT 0.215 2.15 0.42 2.635 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.54 ;
  ANTENNAPARTIALMETALAREA 0.3196 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.3568 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 3.895 2.35 4.835 2.69 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.77 -0.4 13.86 0.4 ;
      RECT 12.43 -0.4 12.77 1.615 ;
      RECT 10.08 -0.4 12.43 0.4 ;
      RECT 9.74 -0.4 10.08 0.575 ;
      RECT 4.725 -0.4 9.74 0.4 ;
      RECT 4.385 -0.4 4.725 0.9 ;
      RECT 1.285 -0.4 4.385 0.4 ;
      RECT 0.945 -0.4 1.285 0.575 ;
      RECT 0 -0.4 0.945 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.775 4.64 13.86 5.44 ;
      RECT 12.435 3.93 12.775 5.44 ;
      RECT 8.935 4.64 12.435 5.44 ;
      RECT 8.595 4.465 8.935 5.44 ;
      RECT 1.2 4.64 8.595 5.44 ;
      RECT 0.86 4.465 1.2 5.44 ;
      RECT 0 4.64 0.86 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 12.635 2.015 12.865 3.595 ;
      RECT 11.645 3.365 12.635 3.595 ;
      RECT 11.415 3.365 11.645 3.945 ;
      RECT 9.395 4.18 11.455 4.41 ;
      RECT 10.455 3.715 11.415 3.945 ;
      RECT 11.14 0.63 11.295 0.86 ;
      RECT 11.14 3.12 11.175 3.46 ;
      RECT 10.91 0.63 11.14 3.46 ;
      RECT 10.9 0.63 10.91 1.04 ;
      RECT 10.835 3.12 10.91 3.46 ;
      RECT 9.495 0.81 10.9 1.04 ;
      RECT 10.455 1.345 10.68 1.77 ;
      RECT 10.45 1.345 10.455 3.945 ;
      RECT 10.225 1.54 10.45 3.945 ;
      RECT 10.115 3.215 10.225 3.555 ;
      RECT 9.73 1.27 9.96 2.875 ;
      RECT 9.035 1.27 9.73 1.5 ;
      RECT 9.68 2.645 9.73 2.875 ;
      RECT 9.45 2.645 9.68 3.555 ;
      RECT 9.265 0.63 9.495 1.04 ;
      RECT 9.165 4.005 9.395 4.41 ;
      RECT 5.88 0.63 9.265 0.86 ;
      RECT 7.855 4.005 9.165 4.235 ;
      RECT 8.805 1.09 9.035 1.5 ;
      RECT 6.67 1.09 8.805 1.32 ;
      RECT 8.57 2.195 8.76 2.535 ;
      RECT 8.34 1.585 8.57 2.535 ;
      RECT 8.315 2.305 8.34 2.535 ;
      RECT 8.085 2.305 8.315 3.77 ;
      RECT 7.85 3.58 7.855 4.235 ;
      RECT 7.625 1.585 7.85 4.235 ;
      RECT 7.62 1.585 7.625 3.81 ;
      RECT 7.175 3.58 7.62 3.81 ;
      RECT 7.16 1.79 7.39 3.35 ;
      RECT 7.13 1.79 7.16 2.02 ;
      RECT 6.795 3.12 7.16 3.35 ;
      RECT 6.9 1.585 7.13 2.02 ;
      RECT 6.67 2.36 6.93 2.7 ;
      RECT 6.685 3.12 6.795 3.78 ;
      RECT 6.565 3.12 6.685 4.41 ;
      RECT 6.44 1.09 6.67 2.89 ;
      RECT 6.455 3.44 6.565 4.41 ;
      RECT 5.255 4.055 6.455 4.41 ;
      RECT 6.175 2.655 6.44 2.89 ;
      RECT 5.3 2.07 6.21 2.42 ;
      RECT 6.075 2.655 6.175 3.425 ;
      RECT 5.945 2.655 6.075 3.48 ;
      RECT 5.765 3.14 5.945 3.48 ;
      RECT 5.65 0.63 5.88 1.75 ;
      RECT 5.735 3.14 5.765 3.825 ;
      RECT 5.535 3.195 5.735 3.825 ;
      RECT 5.54 1.135 5.65 1.75 ;
      RECT 4.155 1.135 5.54 1.365 ;
      RECT 3.44 3.595 5.535 3.825 ;
      RECT 5.07 1.635 5.3 3.365 ;
      RECT 1.66 4.18 5.255 4.41 ;
      RECT 3.695 1.635 5.07 1.865 ;
      RECT 3.9 3.135 5.07 3.365 ;
      RECT 3.925 0.875 4.155 1.365 ;
      RECT 2.45 0.875 3.925 1.105 ;
      RECT 3.67 2.98 3.9 3.365 ;
      RECT 3.465 1.44 3.695 1.865 ;
      RECT 3.21 3.03 3.44 3.825 ;
      RECT 3.18 3.03 3.21 3.26 ;
      RECT 2.95 2.075 3.18 3.26 ;
      RECT 2.75 3.495 2.98 3.95 ;
      RECT 2.91 2.075 2.95 2.305 ;
      RECT 2.68 1.42 2.91 2.305 ;
      RECT 2.125 3.495 2.75 3.725 ;
      RECT 2.45 2.535 2.62 3.265 ;
      RECT 2.39 0.875 2.45 3.265 ;
      RECT 2.22 0.875 2.39 2.765 ;
      RECT 1.99 3.05 2.125 3.725 ;
      RECT 1.895 1.395 1.99 3.725 ;
      RECT 1.76 1.395 1.895 3.28 ;
      RECT 1.505 2.94 1.76 3.28 ;
      RECT 1.43 3.655 1.66 4.41 ;
      RECT 1.38 2.04 1.49 2.38 ;
      RECT 1.235 3.655 1.43 3.885 ;
      RECT 1.235 1.395 1.38 2.38 ;
      RECT 1.15 1.395 1.235 3.885 ;
      RECT 0.52 1.395 1.15 1.625 ;
      RECT 1.005 2.095 1.15 3.885 ;
      RECT 0.18 2.89 1.005 3.23 ;
      RECT 0.18 0.815 0.52 1.625 ;
  END
END CMPR32X1

MACRO CMPR22X1
  CLASS CORE ;
  FOREIGN CMPR22X1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.92 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.8762 ;
  ANTENNAPARTIALMETALAREA 1.1041 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.6481 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.005 1.33 4.235 3.22 ;
      RECT 3.59 1.33 4.005 1.56 ;
      RECT 3.245 2.84 4.005 3.22 ;
      RECT 3.36 1.21 3.59 1.56 ;
      RECT 3.015 2.84 3.245 3.73 ;
     END
  END S

  PIN CO
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.8148 ;
  ANTENNAPARTIALMETALAREA 0.7152 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.5404 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.61 1.845 7.705 2.075 ;
      RECT 7.4 1.38 7.61 2.075 ;
      RECT 7.38 1.38 7.4 3.115 ;
      RECT 7.185 1.845 7.38 3.115 ;
      RECT 7.17 1.845 7.185 3.97 ;
      RECT 6.955 2.885 7.17 3.97 ;
     END
  END CO

  PIN B
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.846 ;
  ANTENNAPARTIALMETALAREA 2.1553 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.8103 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.835 2.52 6.065 3.445 ;
      RECT 5.16 3.215 5.835 3.445 ;
      RECT 4.93 3.215 5.16 4.235 ;
      RECT 2.785 4.005 4.93 4.235 ;
      RECT 3.545 1.8 3.775 2.52 ;
      RECT 2.785 2.29 3.545 2.52 ;
      RECT 2.555 2.29 2.785 4.235 ;
      RECT 2.195 2.29 2.555 2.66 ;
      RECT 2.115 2.29 2.195 2.575 ;
      RECT 1.775 2.235 2.115 2.575 ;
     END
  END B

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.846 ;
  ANTENNAPARTIALMETALAREA 0.2562 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0918 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 4.465 1.82 5.075 2.24 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 7.15 -0.4 7.92 0.4 ;
      RECT 6.92 -0.4 7.15 1.355 ;
      RECT 5.125 -0.4 6.92 0.4 ;
      RECT 6.815 1.125 6.92 1.355 ;
      RECT 6.585 1.125 6.815 1.72 ;
      RECT 4.785 -0.4 5.125 0.575 ;
      RECT 1.36 -0.4 4.785 0.4 ;
      RECT 1.02 -0.4 1.36 0.575 ;
      RECT 0 -0.4 1.02 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 6.48 4.64 7.92 5.44 ;
      RECT 6.14 4.465 6.48 5.44 ;
      RECT 4.78 4.64 6.14 5.44 ;
      RECT 4.44 4.465 4.78 5.44 ;
      RECT 1.28 4.64 4.44 5.44 ;
      RECT 0.94 4.465 1.28 5.44 ;
      RECT 0 4.64 0.94 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 6.525 1.98 6.84 2.32 ;
      RECT 6.35 0.665 6.69 0.895 ;
      RECT 6.35 1.98 6.525 3.905 ;
      RECT 6.295 0.665 6.35 3.905 ;
      RECT 6.12 0.665 6.295 2.21 ;
      RECT 5.625 3.675 6.295 3.905 ;
      RECT 5.6 1.21 5.885 1.55 ;
      RECT 5.395 3.675 5.625 4.085 ;
      RECT 5.545 1.21 5.6 2.985 ;
      RECT 5.37 1.265 5.545 2.985 ;
      RECT 4.7 1.265 5.37 1.495 ;
      RECT 4.7 2.755 5.37 2.985 ;
      RECT 4.47 0.805 4.7 1.495 ;
      RECT 4.47 2.755 4.7 3.775 ;
      RECT 4.365 0.805 4.47 1.035 ;
      RECT 3.68 3.545 4.47 3.775 ;
      RECT 4.025 0.675 4.365 1.035 ;
      RECT 3.13 0.675 4.025 0.905 ;
      RECT 2.9 0.675 3.13 1.955 ;
      RECT 1.385 1.725 2.9 1.955 ;
      RECT 2.44 0.63 2.67 1.035 ;
      RECT 0.925 1.265 2.55 1.495 ;
      RECT 0.465 0.805 2.44 1.035 ;
      RECT 2.095 4.005 2.325 4.405 ;
      RECT 0.465 4.005 2.095 4.235 ;
      RECT 1.5 3.18 1.84 3.52 ;
      RECT 0.925 3.18 1.5 3.41 ;
      RECT 1.155 1.725 1.385 2.56 ;
      RECT 0.695 1.265 0.925 3.41 ;
      RECT 0.235 0.76 0.465 4.235 ;
  END
END CMPR22X1

MACRO BMXX1
  CLASS CORE ;
  FOREIGN BMXX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.54 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN X2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3366 ;
  ANTENNAPARTIALMETALAREA 0.2553 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0759 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.38 2.16 9.84 2.715 ;
     END
  END X2

  PIN S
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3294 ;
  ANTENNAPARTIALMETALAREA 0.2063 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 0.9646 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 6.69 2.185 7.12 2.665 ;
     END
  END S

  PIN PP
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 0.72 ;
  ANTENNAPARTIALMETALAREA 0.6446 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.8726 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 12.305 2.635 12.36 3.635 ;
      RECT 12.075 1.265 12.305 3.635 ;
      RECT 12.02 2.825 12.075 3.635 ;
     END
  END PP

  PIN M1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3006 ;
  ANTENNAPARTIALMETALAREA 0.2544 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0706 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 5.93 1.79 6.46 2.27 ;
     END
  END M1

  PIN M0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3006 ;
  ANTENNAPARTIALMETALAREA 0.2334 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.1236 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 0.8 1.82 1.11 2.54 ;
      RECT 0.77 2.2 0.8 2.54 ;
     END
  END M0

  PIN A
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.3294 ;
  ANTENNAPARTIALMETALAREA 0.221 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 1.0494 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.46 2.01 1.8 2.66 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 12.36 -0.4 12.54 0.4 ;
      RECT 12.02 -0.4 12.36 0.575 ;
      RECT 8.625 -0.4 12.02 0.4 ;
      RECT 8.285 -0.4 8.625 0.575 ;
      RECT 6.605 -0.4 8.285 0.4 ;
      RECT 6.265 -0.4 6.605 0.575 ;
      RECT 1.32 -0.4 6.265 0.4 ;
      RECT 0.98 -0.4 1.32 1.52 ;
      RECT 0 -0.4 0.98 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 11.935 4.64 12.54 5.44 ;
      RECT 11.595 4.465 11.935 5.44 ;
      RECT 9.09 4.64 11.595 5.44 ;
      RECT 6.4 4.465 9.09 5.44 ;
      RECT 1.32 4.64 6.4 5.44 ;
      RECT 0.98 3.92 1.32 5.44 ;
      RECT 0 4.64 0.98 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 11.79 1.085 11.805 2.595 ;
      RECT 11.575 0.665 11.79 2.595 ;
      RECT 11.56 0.665 11.575 1.315 ;
      RECT 11.515 2.365 11.575 2.595 ;
      RECT 10.96 0.665 11.56 0.895 ;
      RECT 11.365 2.365 11.515 3.985 ;
      RECT 11.285 2.365 11.365 4.375 ;
      RECT 11.33 1.65 11.345 2.135 ;
      RECT 11.115 1.125 11.33 2.135 ;
      RECT 11.135 3.755 11.285 4.375 ;
      RECT 9.665 4.145 11.135 4.375 ;
      RECT 11.1 1.125 11.115 1.88 ;
      RECT 10.3 1.125 11.1 1.355 ;
      RECT 10.62 0.63 10.96 0.895 ;
      RECT 10.905 2.855 10.915 3.365 ;
      RECT 10.87 2.855 10.905 3.81 ;
      RECT 10.675 1.585 10.87 3.81 ;
      RECT 10.64 1.585 10.675 3.085 ;
      RECT 8.69 3.58 10.675 3.81 ;
      RECT 10.53 1.585 10.64 1.815 ;
      RECT 9.535 0.63 10.62 0.86 ;
      RECT 10.07 1.125 10.3 3.32 ;
      RECT 9.77 1.46 10.07 1.69 ;
      RECT 9.865 3.09 10.07 3.32 ;
      RECT 9.15 3.06 9.445 3.29 ;
      RECT 9.15 1.43 9.335 1.93 ;
      RECT 5.98 0.805 9.195 1.035 ;
      RECT 9.105 1.43 9.15 3.29 ;
      RECT 8.92 1.7 9.105 3.29 ;
      RECT 8.46 2.995 8.69 3.81 ;
      RECT 8.07 2.995 8.46 3.225 ;
      RECT 7.84 1.265 8.07 3.225 ;
      RECT 7.83 3.695 7.98 3.925 ;
      RECT 7.725 1.265 7.84 1.495 ;
      RECT 7.6 3.695 7.83 4.235 ;
      RECT 5.9 4.005 7.6 4.235 ;
      RECT 7.37 1.725 7.58 3.195 ;
      RECT 7.365 1.725 7.37 3.775 ;
      RECT 7.35 1.265 7.365 3.775 ;
      RECT 7.135 1.265 7.35 1.955 ;
      RECT 7.14 2.965 7.35 3.775 ;
      RECT 5.44 3.545 7.14 3.775 ;
      RECT 7.025 1.265 7.135 1.605 ;
      RECT 5.75 0.63 5.98 1.035 ;
      RECT 5.7 2.83 5.98 3.17 ;
      RECT 5.67 4.005 5.9 4.405 ;
      RECT 5.7 1.33 5.875 1.56 ;
      RECT 4.4 0.63 5.75 0.86 ;
      RECT 5.64 1.33 5.7 3.17 ;
      RECT 3.02 4.175 5.67 4.405 ;
      RECT 5.47 1.33 5.64 3.115 ;
      RECT 5.21 2.21 5.47 2.55 ;
      RECT 5.21 3.545 5.44 3.945 ;
      RECT 4.97 2.85 5.24 3.19 ;
      RECT 3.48 3.715 5.21 3.945 ;
      RECT 4.97 1.09 5.175 1.32 ;
      RECT 4.74 1.09 4.97 3.485 ;
      RECT 3.94 3.255 4.74 3.485 ;
      RECT 4.4 2.795 4.51 3.025 ;
      RECT 4.17 0.63 4.4 3.025 ;
      RECT 3.71 0.63 3.94 3.485 ;
      RECT 2.04 0.63 3.71 0.86 ;
      RECT 3.25 1.09 3.48 3.945 ;
      RECT 3.14 1.09 3.25 1.32 ;
      RECT 2.79 3.03 3.02 4.405 ;
      RECT 2.76 3.03 2.79 3.26 ;
      RECT 2.53 1.09 2.76 3.26 ;
      RECT 2.3 3.49 2.56 3.83 ;
      RECT 2.42 1.09 2.53 1.32 ;
      RECT 2.07 1.55 2.3 3.23 ;
      RECT 2.22 3.46 2.3 3.83 ;
      RECT 2.07 3.46 2.22 3.775 ;
      RECT 2.04 1.55 2.07 1.78 ;
      RECT 1.74 2.89 2.07 3.23 ;
      RECT 0.52 3.46 2.07 3.69 ;
      RECT 1.81 0.63 2.04 1.78 ;
      RECT 1.7 1.035 1.81 1.375 ;
      RECT 0.29 1.455 0.52 3.69 ;
      RECT 0.18 1.455 0.29 1.795 ;
      RECT 0.18 2.83 0.29 3.17 ;
  END
END BMXX1

MACRO BENCX4
  CLASS CORE ;
  FOREIGN BENCX4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 40.26 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN X2
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 5.4561 ;
  ANTENNAPARTIALMETALAREA 2.4333 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.5735 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 27.58 1.345 27.695 1.575 ;
      RECT 27.58 2.625 27.69 2.855 ;
      RECT 27.2 1.345 27.58 2.855 ;
      RECT 23.275 1.345 27.2 1.575 ;
      RECT 23.265 2.625 27.2 2.855 ;
     END
  END X2

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 5.4552 ;
  ANTENNAPARTIALMETALAREA 2.8125 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 12.3967 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 39.975 1.82 40.12 3.22 ;
      RECT 39.97 1.82 39.975 3.24 ;
      RECT 39.74 1.515 39.97 3.24 ;
      RECT 34.95 1.515 39.74 1.745 ;
      RECT 34.94 3.01 39.74 3.24 ;
     END
  END S

  PIN M2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.7776 ;
  ANTENNAPARTIALMETALAREA 3.9836 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 18.603 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.79 4.005 28.985 4.235 ;
      RECT 20.56 4.005 20.79 4.41 ;
      RECT 16.925 4.18 20.56 4.41 ;
      RECT 16.695 4.005 16.925 4.41 ;
      RECT 12.325 4.005 16.695 4.235 ;
      RECT 12.095 4.005 12.325 4.315 ;
     END
  END M2

  PIN M1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 2.0628 ;
  ANTENNAPARTIALMETALAREA 2.583 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.9886 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 16.51 3.43 16.74 3.775 ;
      RECT 12.805 3.545 16.51 3.775 ;
      RECT 12.575 3.075 12.805 3.775 ;
      RECT 9.455 3.105 12.575 3.335 ;
      RECT 9.245 2.94 9.455 3.335 ;
      RECT 9.015 2.56 9.245 3.335 ;
      RECT 7.405 2.965 9.015 3.195 ;
      RECT 7.175 2.58 7.405 3.195 ;
     END
  END M1

  PIN M0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.7532 ;
  ANTENNAPARTIALMETALAREA 2.2095 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.2714 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 13.4 0.635 13.56 1.955 ;
      RECT 13.33 0.635 13.4 2.385 ;
      RECT 12.64 0.635 13.33 0.865 ;
      RECT 13.17 1.725 13.33 2.385 ;
      RECT 12.41 0.635 12.64 1.035 ;
      RECT 10.97 0.805 12.41 1.035 ;
      RECT 10.74 0.805 10.97 2.05 ;
      RECT 8.365 1.82 10.74 2.05 ;
      RECT 8.135 1.82 8.365 2.635 ;
      RECT 8.06 1.955 8.135 2.635 ;
      RECT 7.55 1.955 8.06 2.185 ;
     END
  END M0

  PIN A
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 5.33 ;
  ANTENNAPARTIALMETALAREA 3.3128 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.6159 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.185 1.39 5.085 1.73 ;
      RECT 1.185 2.74 5.085 3.08 ;
      RECT 1.18 1.39 1.185 3.08 ;
      RECT 0.9 1.39 1.18 3.22 ;
      RECT 0.8 1.82 0.9 3.22 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 40.05 -0.4 40.26 0.4 ;
      RECT 39.71 -0.4 40.05 1.11 ;
      RECT 38.69 -0.4 39.71 0.4 ;
      RECT 38.35 -0.4 38.69 1.11 ;
      RECT 37.33 -0.4 38.35 0.4 ;
      RECT 36.99 -0.4 37.33 1.11 ;
      RECT 35.97 -0.4 36.99 0.4 ;
      RECT 35.63 -0.4 35.97 1.11 ;
      RECT 34.61 -0.4 35.63 0.4 ;
      RECT 34.27 -0.4 34.61 1.11 ;
      RECT 33.135 -0.4 34.27 0.4 ;
      RECT 33.135 0.77 33.285 1.11 ;
      RECT 32.795 -0.4 33.135 1.11 ;
      RECT 31.335 -0.4 32.795 0.4 ;
      RECT 32.475 0.77 32.795 1.11 ;
      RECT 30.995 -0.4 31.335 0.575 ;
      RECT 28.375 -0.4 30.995 0.4 ;
      RECT 28.035 -0.4 28.375 0.575 ;
      RECT 27.015 -0.4 28.035 0.4 ;
      RECT 26.675 -0.4 27.015 0.575 ;
      RECT 25.655 -0.4 26.675 0.4 ;
      RECT 25.315 -0.4 25.655 0.575 ;
      RECT 24.295 -0.4 25.315 0.4 ;
      RECT 23.955 -0.4 24.295 0.575 ;
      RECT 22.935 -0.4 23.955 0.4 ;
      RECT 22.595 -0.4 22.935 0.575 ;
      RECT 21.575 -0.4 22.595 0.4 ;
      RECT 21.235 -0.4 21.575 0.575 ;
      RECT 15.895 -0.4 21.235 0.4 ;
      RECT 15.605 -0.4 15.895 0.575 ;
      RECT 15.605 0.98 15.895 1.32 ;
      RECT 15.375 -0.4 15.605 1.32 ;
      RECT 15.085 -0.4 15.375 0.575 ;
      RECT 15.085 0.98 15.375 1.32 ;
      RECT 12.18 -0.4 15.085 0.4 ;
      RECT 11.84 -0.4 12.18 0.575 ;
      RECT 8.84 -0.4 11.84 0.4 ;
      RECT 8.5 -0.4 8.84 0.575 ;
      RECT 7.225 -0.4 8.5 0.4 ;
      RECT 6.885 -0.4 7.225 0.95 ;
      RECT 5.725 -0.4 6.885 0.4 ;
      RECT 5.385 -0.4 5.725 0.95 ;
      RECT 4.445 -0.4 5.385 0.4 ;
      RECT 4.105 -0.4 4.445 0.95 ;
      RECT 3.165 -0.4 4.105 0.4 ;
      RECT 2.825 -0.4 3.165 0.95 ;
      RECT 1.88 -0.4 2.825 0.4 ;
      RECT 1.54 -0.4 1.88 0.95 ;
      RECT 0.6 -0.4 1.54 0.4 ;
      RECT 0.26 -0.4 0.6 0.95 ;
      RECT 0 -0.4 0.26 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 40.045 4.64 40.26 5.44 ;
      RECT 39.705 3.775 40.045 5.44 ;
      RECT 38.685 4.64 39.705 5.44 ;
      RECT 38.345 3.775 38.685 5.44 ;
      RECT 37.325 4.64 38.345 5.44 ;
      RECT 36.985 3.775 37.325 5.44 ;
      RECT 35.965 4.64 36.985 5.44 ;
      RECT 35.625 3.775 35.965 5.44 ;
      RECT 34.6 4.64 35.625 5.44 ;
      RECT 34.26 3.775 34.6 5.44 ;
      RECT 33.24 4.64 34.26 5.44 ;
      RECT 32.9 3.825 33.24 5.44 ;
      RECT 30.285 4.64 32.9 5.44 ;
      RECT 29.945 3.825 30.285 5.44 ;
      RECT 28.37 4.64 29.945 5.44 ;
      RECT 28.03 4.465 28.37 5.44 ;
      RECT 27.01 4.64 28.03 5.44 ;
      RECT 26.67 4.465 27.01 5.44 ;
      RECT 25.65 4.64 26.67 5.44 ;
      RECT 25.31 4.465 25.65 5.44 ;
      RECT 24.29 4.64 25.31 5.44 ;
      RECT 23.95 4.465 24.29 5.44 ;
      RECT 22.925 4.64 23.95 5.44 ;
      RECT 22.585 4.465 22.925 5.44 ;
      RECT 21.565 4.64 22.585 5.44 ;
      RECT 21.225 4.465 21.565 5.44 ;
      RECT 16.465 4.64 21.225 5.44 ;
      RECT 16.125 4.465 16.465 5.44 ;
      RECT 14.855 4.64 16.125 5.44 ;
      RECT 14.515 4.465 14.855 5.44 ;
      RECT 13.23 4.64 14.515 5.44 ;
      RECT 12.89 4.465 13.23 5.44 ;
      RECT 11.515 4.64 12.89 5.44 ;
      RECT 11.285 4.005 11.515 5.44 ;
      RECT 9.71 4.64 11.285 5.44 ;
      RECT 9.37 4.465 9.71 5.44 ;
      RECT 7.06 4.64 9.37 5.44 ;
      RECT 6.72 4.465 7.06 5.44 ;
      RECT 5.725 4.64 6.72 5.44 ;
      RECT 5.385 3.85 5.725 5.44 ;
      RECT 4.445 4.64 5.385 5.44 ;
      RECT 4.105 3.85 4.445 5.44 ;
      RECT 3.165 4.64 4.105 5.44 ;
      RECT 2.825 3.85 3.165 5.44 ;
      RECT 1.88 4.64 2.825 5.44 ;
      RECT 1.54 3.85 1.88 5.44 ;
      RECT 0.6 4.64 1.54 5.44 ;
      RECT 0.26 3.85 0.6 5.44 ;
      RECT 0 4.64 0.26 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 34.5 2.06 38.605 2.29 ;
      RECT 34.415 1.515 34.5 2.29 ;
      RECT 34.27 1.515 34.415 3.025 ;
      RECT 33.59 1.515 34.27 1.745 ;
      RECT 34.185 2.06 34.27 3.025 ;
      RECT 33.58 2.795 34.185 3.025 ;
      RECT 33.36 2.19 33.84 2.42 ;
      RECT 33.35 1.35 33.36 2.42 ;
      RECT 33.13 1.35 33.35 3.595 ;
      RECT 29.355 1.35 33.13 1.58 ;
      RECT 33.12 2.19 33.13 3.595 ;
      RECT 31.55 3.365 33.12 3.595 ;
      RECT 32.66 1.99 32.89 2.855 ;
      RECT 30.895 2.625 32.66 2.855 ;
      RECT 30.415 0.805 32.095 1.035 ;
      RECT 31.32 3.12 31.55 4.405 ;
      RECT 29.47 3.365 31.32 3.595 ;
      RECT 30.665 1.81 30.895 3.11 ;
      RECT 28.7 1.81 30.665 2.04 ;
      RECT 29.01 2.88 30.665 3.11 ;
      RECT 28.55 2.27 30.435 2.5 ;
      RECT 30.185 0.63 30.415 1.035 ;
      RECT 29.095 0.63 30.185 0.86 ;
      RECT 29.24 3.365 29.47 4.225 ;
      RECT 28.78 2.88 29.01 3.775 ;
      RECT 20.3 3.545 28.78 3.775 ;
      RECT 28.47 0.805 28.7 2.04 ;
      RECT 28.32 2.27 28.55 3.315 ;
      RECT 21.005 0.805 28.47 1.035 ;
      RECT 21.015 3.085 28.32 3.315 ;
      RECT 22.3 1.89 26.93 2.12 ;
      RECT 22.2 1.89 22.3 2.855 ;
      RECT 22.07 1.29 22.2 2.855 ;
      RECT 21.97 1.29 22.07 2.12 ;
      RECT 21.905 2.625 22.07 2.855 ;
      RECT 20.545 1.89 21.73 2.12 ;
      RECT 20.785 2.535 21.015 3.315 ;
      RECT 20.775 0.63 21.005 1.035 ;
      RECT 20.135 2.535 20.785 2.765 ;
      RECT 16.42 0.63 20.775 0.86 ;
      RECT 20.315 1.09 20.545 2.305 ;
      RECT 17.425 1.09 20.315 1.32 ;
      RECT 19.695 2.075 20.315 2.305 ;
      RECT 20.07 3.545 20.3 3.95 ;
      RECT 19.235 1.55 20.085 1.78 ;
      RECT 17.395 3.72 20.07 3.95 ;
      RECT 19.465 2.075 19.695 3.49 ;
      RECT 17.705 3.26 19.465 3.49 ;
      RECT 19.005 1.55 19.235 3.03 ;
      RECT 17.145 1.55 19.005 1.78 ;
      RECT 17.395 2.8 19.005 3.03 ;
      RECT 16.935 2.27 18.775 2.5 ;
      RECT 17.165 2.8 17.395 3.2 ;
      RECT 17.165 3.49 17.395 3.95 ;
      RECT 16.285 2.97 17.165 3.2 ;
      RECT 16.985 3.49 17.165 3.72 ;
      RECT 16.915 1.265 17.145 1.78 ;
      RECT 16.705 2.27 16.935 2.74 ;
      RECT 16.705 1.265 16.915 1.495 ;
      RECT 14.66 2.51 16.705 2.74 ;
      RECT 16.19 0.63 16.42 2.215 ;
      RECT 16.055 2.97 16.285 3.26 ;
      RECT 14.51 1.985 16.19 2.215 ;
      RECT 15.365 3.03 16.055 3.26 ;
      RECT 14.43 2.51 14.66 3.315 ;
      RECT 14.28 0.715 14.51 2.215 ;
      RECT 13.265 3.085 14.43 3.315 ;
      RECT 14.125 1.985 14.28 2.215 ;
      RECT 13.895 1.985 14.125 2.855 ;
      RECT 13.69 2.625 13.895 2.855 ;
      RECT 13.035 2.615 13.265 3.315 ;
      RECT 12.935 1.095 13.1 1.495 ;
      RECT 12.935 2.615 13.035 2.845 ;
      RECT 12.87 1.095 12.935 2.845 ;
      RECT 12.705 1.265 12.87 2.845 ;
      RECT 11.99 2.545 12.705 2.775 ;
      RECT 11.515 1.265 11.77 1.495 ;
      RECT 11.285 1.265 11.515 2.51 ;
      RECT 11.015 2.28 11.285 2.51 ;
      RECT 10.665 2.28 11.015 2.87 ;
      RECT 9.63 2.28 10.665 2.51 ;
      RECT 9.34 0.635 10.48 0.865 ;
      RECT 6.83 1.355 10.48 1.585 ;
      RECT 8.335 3.565 10.47 3.795 ;
      RECT 9.11 0.635 9.34 1.035 ;
      RECT 7.74 0.805 9.11 1.035 ;
      RECT 8.105 3.5 8.335 4.31 ;
      RECT 6.83 3.5 8.105 3.73 ;
      RECT 6.6 1.355 6.83 3.73 ;
      RECT 6.26 2.09 6.6 2.43 ;
      RECT 6.03 1.39 6.37 1.73 ;
      RECT 6.03 2.74 6.37 3.08 ;
      RECT 6.025 1.5 6.03 1.73 ;
      RECT 6.025 2.74 6.03 2.97 ;
      RECT 5.795 1.5 6.025 2.97 ;
      RECT 5.325 2.155 5.795 2.385 ;
      RECT 4.515 2.1 5.325 2.44 ;
      RECT 3.12 2.155 4.515 2.385 ;
      RECT 2.31 2.1 3.12 2.44 ;
  END
END BENCX4

MACRO BENCX2
  CLASS CORE ;
  FOREIGN BENCX2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 27.06 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BENCX4 ;

  PIN X2
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.1688 ;
  ANTENNAPARTIALMETALAREA 1.2378 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 5.6551 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 17.945 1.265 18.855 1.495 ;
      RECT 17.945 2.625 18.285 2.855 ;
      RECT 17.715 1.265 17.945 2.855 ;
      RECT 16.985 1.265 17.715 1.495 ;
      RECT 17.605 2.38 17.715 2.855 ;
      RECT 17.02 2.625 17.605 2.855 ;
      RECT 16.64 2.38 17.02 2.855 ;
      RECT 16.425 2.625 16.64 2.855 ;
     END
  END X2

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.2076 ;
  ANTENNAPARTIALMETALAREA 1.7563 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.4836 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 26.11 2.965 26.185 3.195 ;
      RECT 25.96 1.315 26.11 3.195 ;
      RECT 25.955 1.315 25.96 3.72 ;
      RECT 25.88 1.26 25.955 3.72 ;
      RECT 25.72 1.26 25.88 1.545 ;
      RECT 25.62 2.965 25.88 3.72 ;
      RECT 25.38 1.205 25.72 1.545 ;
      RECT 25.525 2.965 25.62 3.22 ;
      RECT 24.635 2.965 25.525 3.195 ;
      RECT 24.28 1.26 25.38 1.545 ;
      RECT 24.52 2.965 24.635 3.22 ;
      RECT 24.29 2.965 24.52 3.74 ;
      RECT 24.18 3.4 24.29 3.74 ;
      RECT 23.94 1.205 24.28 1.545 ;
     END
  END S

  PIN M2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.4212 ;
  ANTENNAPARTIALMETALAREA 2.5104 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 11.8137 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 19.545 4.055 19.655 4.285 ;
      RECT 19.315 4.005 19.545 4.285 ;
      RECT 15.135 4.005 19.315 4.235 ;
      RECT 14.905 4.005 15.135 4.41 ;
      RECT 11.14 4.18 14.905 4.41 ;
      RECT 10.91 4.005 11.14 4.41 ;
      RECT 9.685 4.005 10.91 4.235 ;
      RECT 9.455 4.005 9.685 4.315 ;
      RECT 9.22 4.005 9.455 4.235 ;
     END
  END M2

  PIN M1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.1088 ;
  ANTENNAPARTIALMETALAREA 2.1068 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.9534 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 10.72 2.77 11.775 3 ;
      RECT 10.49 2.77 10.72 3.775 ;
      RECT 8.325 3.545 10.49 3.775 ;
      RECT 8.095 3.545 8.325 4.36 ;
      RECT 5.8 3.545 8.095 3.775 ;
      RECT 5.8 2.305 6.08 2.535 ;
      RECT 5.57 2.305 5.8 3.775 ;
      RECT 5.495 2.965 5.57 3.195 ;
     END
  END M1

  PIN M0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 1.017 ;
  ANTENNAPARTIALMETALAREA 1.7384 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.0136 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 8.895 0.63 10.07 0.86 ;
      RECT 8.665 0.63 8.895 1.035 ;
      RECT 7.78 0.805 8.665 1.035 ;
      RECT 7.57 0.805 7.78 1.285 ;
      RECT 7.34 0.805 7.57 2.235 ;
      RECT 6.54 2.005 7.34 2.235 ;
      RECT 6.31 1.845 6.54 2.235 ;
      RECT 5.14 1.845 6.31 2.075 ;
      RECT 4.91 1.845 5.14 2.635 ;
      RECT 4.835 2.405 4.91 2.635 ;
     END
  END M0

  PIN A
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 3.2076 ;
  ANTENNAPARTIALMETALAREA 2.1871 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 8.0454 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 2.35 0.835 2.69 1.645 ;
      RECT 2.35 3.09 2.69 3.955 ;
      RECT 1.25 1.415 2.35 1.645 ;
      RECT 1.535 3.09 2.35 3.32 ;
      RECT 1.25 2.94 1.535 3.32 ;
      RECT 0.91 0.835 1.25 3.955 ;
      RECT 0.875 2.405 0.91 2.635 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 26.385 -0.4 27.06 0.4 ;
      RECT 26.155 -0.4 26.385 0.955 ;
      RECT 25 -0.4 26.155 0.4 ;
      RECT 24.66 -0.4 25 0.965 ;
      RECT 23.52 -0.4 24.66 0.4 ;
      RECT 23.18 -0.4 23.52 0.575 ;
      RECT 22.4 -0.4 23.18 0.4 ;
      RECT 22.06 -0.4 22.4 0.575 ;
      RECT 20.875 -0.4 22.06 0.4 ;
      RECT 20.535 -0.4 20.875 0.575 ;
      RECT 18.09 -0.4 20.535 0.4 ;
      RECT 17.75 -0.4 18.09 0.575 ;
      RECT 16.565 -0.4 17.75 0.4 ;
      RECT 16.225 -0.4 16.565 0.575 ;
      RECT 11.91 -0.4 16.225 0.4 ;
      RECT 11.57 -0.4 11.91 0.575 ;
      RECT 10.53 -0.4 11.57 0.4 ;
      RECT 10.3 -0.4 10.53 1.38 ;
      RECT 8.43 -0.4 10.3 0.4 ;
      RECT 10.05 1.15 10.3 1.38 ;
      RECT 8.09 -0.4 8.43 0.575 ;
      RECT 4.97 -0.4 8.09 0.4 ;
      RECT 4.63 -0.4 4.97 0.575 ;
      RECT 3.45 -0.4 4.63 0.4 ;
      RECT 3.11 -0.4 3.45 1.09 ;
      RECT 1.97 -0.4 3.11 0.4 ;
      RECT 1.63 -0.4 1.97 1.05 ;
      RECT 0.53 -0.4 1.63 0.4 ;
      RECT 0.19 -0.4 0.53 1.49 ;
      RECT 0 -0.4 0.19 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 26.625 4.64 27.06 5.44 ;
      RECT 26.395 3.55 26.625 5.44 ;
      RECT 25.24 4.64 26.395 5.44 ;
      RECT 24.9 3.55 25.24 5.44 ;
      RECT 23.76 4.64 24.9 5.44 ;
      RECT 23.42 3.43 23.76 5.44 ;
      RECT 22.16 4.64 23.42 5.44 ;
      RECT 21.82 4.465 22.16 5.44 ;
      RECT 20.28 4.64 21.82 5.44 ;
      RECT 19.94 4.465 20.28 5.44 ;
      RECT 19.085 4.64 19.94 5.44 ;
      RECT 18.745 4.465 19.085 5.44 ;
      RECT 17.525 4.64 18.745 5.44 ;
      RECT 17.185 4.465 17.525 5.44 ;
      RECT 16.005 4.64 17.185 5.44 ;
      RECT 15.665 4.465 16.005 5.44 ;
      RECT 10.68 4.64 15.665 5.44 ;
      RECT 10.34 4.465 10.68 5.44 ;
      RECT 7.795 4.64 10.34 5.44 ;
      RECT 7.565 4.005 7.795 5.44 ;
      RECT 6.29 4.64 7.565 5.44 ;
      RECT 5.95 4.465 6.29 5.44 ;
      RECT 4.93 4.64 5.95 5.44 ;
      RECT 4.59 4.465 4.93 5.44 ;
      RECT 3.41 4.64 4.59 5.44 ;
      RECT 3.07 4.02 3.41 5.44 ;
      RECT 1.97 4.64 3.07 5.44 ;
      RECT 1.63 3.55 1.97 5.44 ;
      RECT 0.53 4.64 1.63 5.44 ;
      RECT 0.19 3.55 0.53 5.44 ;
      RECT 0 4.64 0.19 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 24.04 2.1 24.85 2.44 ;
      RECT 23.295 2.155 24.04 2.385 ;
      RECT 23.065 1.285 23.295 3.025 ;
      RECT 22.62 1.285 23.065 1.515 ;
      RECT 22.58 2.795 23.065 3.025 ;
      RECT 22.215 2.065 22.555 2.405 ;
      RECT 21.69 2.12 22.215 2.35 ;
      RECT 21.46 1.445 21.69 3.615 ;
      RECT 21.41 0.985 21.635 1.215 ;
      RECT 20.885 1.445 21.46 1.675 ;
      RECT 19.665 3.385 21.46 3.615 ;
      RECT 21.18 0.805 21.41 1.215 ;
      RECT 20.34 2.36 21.23 2.59 ;
      RECT 20.26 0.805 21.18 1.035 ;
      RECT 20.655 1.35 20.885 1.675 ;
      RECT 19.565 1.35 20.655 1.58 ;
      RECT 20.11 1.81 20.34 3.11 ;
      RECT 20.03 0.63 20.26 1.035 ;
      RECT 19.33 1.81 20.11 2.04 ;
      RECT 19.205 2.88 20.11 3.11 ;
      RECT 19.575 0.63 20.03 0.86 ;
      RECT 18.745 2.3 19.88 2.53 ;
      RECT 19.435 3.385 19.665 3.775 ;
      RECT 19.1 0.805 19.33 2.04 ;
      RECT 18.975 2.88 19.205 3.775 ;
      RECT 15.675 0.805 19.1 1.035 ;
      RECT 14.67 3.545 18.975 3.775 ;
      RECT 18.515 2.3 18.745 3.315 ;
      RECT 14.67 3.085 18.515 3.315 ;
      RECT 15.745 1.89 16.71 2.12 ;
      RECT 15.515 1.29 15.745 2.12 ;
      RECT 15.445 0.63 15.675 1.035 ;
      RECT 15.46 1.89 15.515 2.12 ;
      RECT 15.23 1.89 15.46 2.855 ;
      RECT 12.81 0.63 15.445 0.86 ;
      RECT 14.905 2.625 15.23 2.855 ;
      RECT 14.21 1.09 14.72 1.32 ;
      RECT 14.44 2.545 14.67 3.315 ;
      RECT 14.44 3.545 14.67 3.945 ;
      RECT 11.805 3.715 14.44 3.945 ;
      RECT 13.98 1.09 14.21 3.485 ;
      RECT 13.09 1.09 13.98 1.32 ;
      RECT 12.525 3.255 13.98 3.485 ;
      RECT 13.52 1.64 13.75 3.025 ;
      RECT 12.86 1.64 13.52 1.87 ;
      RECT 12.295 2.795 13.52 3.025 ;
      RECT 12.695 2.265 13.29 2.495 ;
      RECT 12.63 1.265 12.86 1.87 ;
      RECT 12.58 0.63 12.81 1.035 ;
      RECT 12.465 2.265 12.695 2.54 ;
      RECT 12.37 1.265 12.63 1.495 ;
      RECT 11.735 0.805 12.58 1.035 ;
      RECT 10.26 2.31 12.465 2.54 ;
      RECT 12.065 2.795 12.295 3.46 ;
      RECT 11.735 1.715 12.065 1.945 ;
      RECT 11.185 3.23 12.065 3.46 ;
      RECT 11.505 0.805 11.735 1.945 ;
      RECT 11.095 1.715 11.505 1.945 ;
      RECT 10.955 3.23 11.185 3.655 ;
      RECT 10.865 0.95 11.095 1.945 ;
      RECT 9.76 1.715 10.865 1.945 ;
      RECT 10.03 2.31 10.26 3.315 ;
      RECT 8.775 3.085 10.03 3.315 ;
      RECT 9.53 1.715 9.76 2.855 ;
      RECT 9.355 1.15 9.675 1.38 ;
      RECT 9.255 2.625 9.53 2.855 ;
      RECT 9.125 1.15 9.355 1.495 ;
      RECT 8.775 1.265 9.125 1.495 ;
      RECT 8.545 1.265 8.775 3.315 ;
      RECT 8.27 3.085 8.545 3.315 ;
      RECT 8.025 1.535 8.255 2.7 ;
      RECT 7.445 2.47 8.025 2.7 ;
      RECT 7.215 2.47 7.445 3.225 ;
      RECT 7.165 2.995 7.215 3.225 ;
      RECT 6.8 2.995 7.165 3.315 ;
      RECT 7 1.545 7.11 1.775 ;
      RECT 6.945 0.825 7.09 1.055 ;
      RECT 4.97 4.005 7.05 4.235 ;
      RECT 6.77 1.385 7 1.775 ;
      RECT 6.715 0.825 6.945 1.155 ;
      RECT 6.28 2.995 6.8 3.225 ;
      RECT 4.67 1.385 6.77 1.615 ;
      RECT 5.39 0.925 6.715 1.155 ;
      RECT 4.74 3.025 4.97 4.235 ;
      RECT 3.895 3.025 4.74 3.255 ;
      RECT 4.44 1.385 4.67 2.01 ;
      RECT 3.895 1.78 4.44 2.01 ;
      RECT 4.06 0.845 4.21 1.185 ;
      RECT 3.79 3.55 4.13 4.36 ;
      RECT 3.83 0.845 4.06 1.55 ;
      RECT 3.665 1.78 3.895 3.255 ;
      RECT 3.155 1.32 3.83 1.55 ;
      RECT 3.155 3.55 3.79 3.78 ;
      RECT 3.555 1.78 3.665 2.12 ;
      RECT 2.925 1.32 3.155 3.78 ;
      RECT 2.115 2.1 2.925 2.44 ;
  END
END BENCX2

MACRO BENCX1
  CLASS CORE ;
  FOREIGN BENCX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 20.46 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;
  LEQ BENCX4 ;

  PIN X2
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.6633 ;
  ANTENNAPARTIALMETALAREA 0.6617 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 2.9839 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 14.06 1.265 14.29 2.855 ;
      RECT 13.785 1.265 14.06 1.495 ;
      RECT 13.9 2.38 14.06 2.855 ;
      RECT 13.34 2.38 13.9 2.66 ;
     END
  END X2

  PIN S
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.566 ;
  ANTENNAPARTIALMETALAREA 0.9853 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 4.6322 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 20.015 1.315 20.245 3.22 ;
      RECT 19.545 1.315 20.015 1.545 ;
      RECT 19.56 2.99 20.015 3.22 ;
      RECT 19.33 2.99 19.56 3.74 ;
      RECT 19.205 1.205 19.545 1.545 ;
      RECT 19.28 3.22 19.33 3.74 ;
      RECT 19.22 3.4 19.28 3.74 ;
     END
  END S

  PIN M2
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.2862 ;
  ANTENNAPARTIALMETALAREA 2.2069 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 10.3774 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 15.67 4.055 15.915 4.285 ;
      RECT 15.44 4.055 15.67 4.35 ;
      RECT 14.075 4.12 15.44 4.35 ;
      RECT 13.94 4.06 14.075 4.35 ;
      RECT 13.71 4.005 13.94 4.35 ;
      RECT 12.8 4.005 13.71 4.235 ;
      RECT 12.57 4.005 12.8 4.41 ;
      RECT 9.715 4.18 12.57 4.41 ;
      RECT 9.485 4.005 9.715 4.41 ;
      RECT 7.705 4.005 9.485 4.235 ;
      RECT 7.475 4.005 7.705 4.315 ;
      RECT 6.965 4.005 7.475 4.235 ;
     END
  END M2

  PIN M1
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5526 ;
  ANTENNAPARTIALMETALAREA 1.9815 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 9.0418 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 9.07 2.77 10.115 3 ;
      RECT 8.84 2.77 9.07 3.775 ;
      RECT 6.635 3.545 8.84 3.775 ;
      RECT 6.295 3.545 6.635 3.83 ;
      RECT 4.315 3.545 6.295 3.775 ;
      RECT 4.085 2.75 4.315 3.775 ;
      RECT 3.905 2.75 4.085 3.22 ;
      RECT 3.44 2.94 3.905 3.22 ;
     END
  END M1

  PIN M0
  DIRECTION INPUT ;
  ANTENNAGATEAREA 0.5526 ;
  ANTENNAPARTIALMETALAREA 1.4858 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 7.0914 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 7.25 0.785 7.695 1.015 ;
      RECT 7.02 0.785 7.25 1.035 ;
      RECT 5.62 0.805 7.02 1.035 ;
      RECT 5.39 0.805 5.62 2.455 ;
      RECT 3.215 2.225 5.39 2.455 ;
      RECT 2.985 2.225 3.215 2.635 ;
      RECT 2.855 2.405 2.985 2.635 ;
     END
  END M0

  PIN A
  DIRECTION OUTPUT ;
  ANTENNADIFFAREA 1.286 ;
  ANTENNAPARTIALMETALAREA 0.7159 LAYER Metal1 ;
  ANTENNAPARTIALMETALSIDEAREA 3.4079 LAYER Metal1 ;
     PORT
      LAYER Metal1 ;
      RECT 1.145 2.74 1.2 3.08 ;
      RECT 0.82 1.46 1.16 1.8 ;
      RECT 0.875 2.74 1.145 3.195 ;
      RECT 0.86 2.74 0.875 3.08 ;
      RECT 0.555 2.74 0.86 2.97 ;
      RECT 0.8 1.54 0.82 1.8 ;
      RECT 0.555 1.57 0.8 1.8 ;
      RECT 0.325 1.57 0.555 2.97 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.265 -0.4 20.46 0.4 ;
      RECT 19.925 -0.4 20.265 0.965 ;
      RECT 18.785 -0.4 19.925 0.4 ;
      RECT 18.445 -0.4 18.785 0.575 ;
      RECT 17.625 -0.4 18.445 0.4 ;
      RECT 17.285 -0.4 17.625 0.575 ;
      RECT 16.335 -0.4 17.285 0.4 ;
      RECT 15.995 -0.4 16.335 0.575 ;
      RECT 14.885 -0.4 15.995 0.4 ;
      RECT 14.545 -0.4 14.885 0.575 ;
      RECT 13.365 -0.4 14.545 0.4 ;
      RECT 13.025 -0.4 13.365 0.575 ;
      RECT 9.005 -0.4 13.025 0.4 ;
      RECT 8.665 -0.4 9.005 0.575 ;
      RECT 6.735 -0.4 8.665 0.4 ;
      RECT 6.395 -0.4 6.735 0.575 ;
      RECT 4.66 -0.4 6.395 0.4 ;
      RECT 4.32 -0.4 4.66 0.575 ;
      RECT 3.14 -0.4 4.32 0.4 ;
      RECT 2.8 -0.4 3.14 0.575 ;
      RECT 1.84 -0.4 2.8 0.4 ;
      RECT 1.5 -0.4 1.84 0.575 ;
      RECT 0.52 -0.4 1.5 0.4 ;
      RECT 0.18 -0.4 0.52 1.05 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 20.28 4.64 20.46 5.44 ;
      RECT 19.94 3.595 20.28 5.44 ;
      RECT 18.8 4.64 19.94 5.44 ;
      RECT 18.46 4.465 18.8 5.44 ;
      RECT 16.485 4.64 18.46 5.44 ;
      RECT 16.145 4.465 16.485 5.44 ;
      RECT 13.48 4.64 16.145 5.44 ;
      RECT 13.14 4.465 13.48 5.44 ;
      RECT 8.915 4.64 13.14 5.44 ;
      RECT 8.575 4.465 8.915 5.44 ;
      RECT 6.065 4.64 8.575 5.44 ;
      RECT 5.835 4.005 6.065 5.44 ;
      RECT 4.465 4.64 5.835 5.44 ;
      RECT 4.125 4.465 4.465 5.44 ;
      RECT 1.88 4.64 4.125 5.44 ;
      RECT 1.54 4.465 1.88 5.44 ;
      RECT 0.52 4.64 1.54 5.44 ;
      RECT 0.18 3.47 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
  OBS
      LAYER Metal1 ;
      RECT 18.965 2.1 19.305 2.44 ;
      RECT 18.335 2.155 18.965 2.385 ;
      RECT 18.105 1.21 18.335 3.225 ;
      RECT 17.885 1.21 18.105 1.44 ;
      RECT 17.805 2.995 18.105 3.225 ;
      RECT 17.575 2.1 17.875 2.44 ;
      RECT 17.55 1.6 17.575 3.69 ;
      RECT 17.345 1.6 17.55 3.98 ;
      RECT 15.765 1.6 17.345 1.83 ;
      RECT 17.32 3.46 17.345 3.98 ;
      RECT 15.67 3.46 17.32 3.69 ;
      RECT 16.255 2.06 17.115 2.29 ;
      RECT 16.29 1.14 16.965 1.37 ;
      RECT 16.06 0.805 16.29 1.37 ;
      RECT 16.025 2.06 16.255 3.215 ;
      RECT 15.76 0.805 16.06 1.035 ;
      RECT 14.755 2.06 16.025 2.29 ;
      RECT 15.21 2.985 16.025 3.215 ;
      RECT 14.75 2.525 15.795 2.755 ;
      RECT 15.535 1.35 15.765 1.83 ;
      RECT 15.53 0.63 15.76 1.035 ;
      RECT 15.44 3.46 15.67 3.81 ;
      RECT 15.265 1.35 15.535 1.58 ;
      RECT 15.245 0.63 15.53 0.86 ;
      RECT 14.98 2.985 15.21 3.775 ;
      RECT 12.34 3.545 14.98 3.775 ;
      RECT 14.525 0.805 14.755 2.29 ;
      RECT 14.52 2.525 14.75 3.315 ;
      RECT 12.8 0.805 14.525 1.035 ;
      RECT 12.34 3.085 14.52 3.315 ;
      RECT 12.805 1.89 13.83 2.12 ;
      RECT 12.805 2.625 12.915 2.855 ;
      RECT 12.575 1.89 12.805 2.855 ;
      RECT 12.57 0.63 12.8 1.035 ;
      RECT 12.34 1.89 12.575 2.12 ;
      RECT 11.085 0.63 12.57 0.86 ;
      RECT 12.11 1.115 12.34 2.12 ;
      RECT 12.11 2.525 12.34 3.315 ;
      RECT 12.11 3.545 12.34 3.945 ;
      RECT 9.945 3.715 12.11 3.945 ;
      RECT 11.65 1.09 11.88 3.485 ;
      RECT 11.5 1.09 11.65 1.405 ;
      RECT 10.805 3.255 11.65 3.485 ;
      RECT 9.985 1.175 11.5 1.405 ;
      RECT 11.19 1.64 11.42 3.025 ;
      RECT 9.67 1.64 11.19 1.87 ;
      RECT 10.575 2.795 11.19 3.025 ;
      RECT 10.73 0.63 11.085 0.945 ;
      RECT 9.72 2.1 10.88 2.33 ;
      RECT 9.465 0.715 10.73 0.945 ;
      RECT 10.345 2.795 10.575 3.46 ;
      RECT 9.53 3.23 10.345 3.46 ;
      RECT 9.49 2.1 9.72 2.54 ;
      RECT 9.44 1.32 9.67 1.87 ;
      RECT 9.3 3.23 9.53 3.655 ;
      RECT 8.61 2.31 9.49 2.54 ;
      RECT 9.235 0.715 9.465 1.035 ;
      RECT 9.225 1.32 9.44 1.55 ;
      RECT 8.985 0.805 9.235 1.035 ;
      RECT 8.985 1.85 9.205 2.08 ;
      RECT 8.755 0.805 8.985 2.08 ;
      RECT 8.295 1.85 8.755 2.08 ;
      RECT 8.38 2.31 8.61 3.315 ;
      RECT 7.58 3.085 8.38 3.315 ;
      RECT 8.15 1.315 8.295 2.08 ;
      RECT 8.065 1.315 8.15 2.855 ;
      RECT 7.905 1.315 8.065 1.545 ;
      RECT 7.92 1.85 8.065 2.855 ;
      RECT 7.81 2.625 7.92 2.855 ;
      RECT 7.35 1.315 7.58 3.315 ;
      RECT 7.205 1.315 7.35 1.545 ;
      RECT 6.525 3.06 7.35 3.29 ;
      RECT 5.85 1.27 6.08 3.28 ;
      RECT 4.645 3.05 5.85 3.28 ;
      RECT 3.34 4.005 5.265 4.235 ;
      RECT 2.5 1.765 5.16 1.995 ;
      RECT 4.875 0.805 5.105 1.33 ;
      RECT 3.56 0.805 4.875 1.035 ;
      RECT 3.205 3.45 3.34 4.235 ;
      RECT 3.11 3.06 3.205 4.235 ;
      RECT 2.975 3.06 3.11 3.68 ;
      RECT 2.5 3.06 2.975 3.29 ;
      RECT 1.67 3.525 2.64 3.755 ;
      RECT 1.67 1.305 2.6 1.535 ;
      RECT 2.27 1.765 2.5 3.29 ;
      RECT 1.93 2.1 2.27 2.44 ;
      RECT 1.44 1.305 1.67 3.755 ;
      RECT 0.79 2.1 1.44 2.44 ;
  END
END BENCX1


MACRO PCORNERDG
    CLASS ENDCAP BOTTOMLEFT ;
    FOREIGN PCORNERDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 235.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE corner ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 235.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 235.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 235.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 235.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 235.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 235.000 235.000 ;
    END
END PCORNERDG

MACRO PDIDGZ
    CLASS PAD ;
    FOREIGN PDIDGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INPUT ;
	AntennaGateArea 6.000000 ;
	AntennaDiffArea 2502.650200 ;
        PORT
        LAYER Metal1 ;
        RECT  18.550 0.000 22.460 1.580 ;
        LAYER Metal2 ;
        RECT  18.550 0.000 22.460 1.580 ;
        END
    END PAD
    PIN C
        DIRECTION OUTPUT ;
	AntennaDiffArea 16.200000 ;
        PORT
        LAYER Metal1 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal2 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal3 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal4 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal5 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal6 ;
        RECT  32.170 234.400 34.170 235.000 ;
        END
    END C
    OBS
        LAYER Metal1 ;
        RECT  34.400 0.000 40.000 235.000 ;
        RECT  31.940 0.000 34.400 234.170 ;
        RECT  22.690 0.000 31.940 235.000 ;
        RECT  18.320 1.810 22.690 235.000 ;
        RECT  0.000 0.000 18.320 235.000 ;
        LAYER Via12 ;
        RECT  32.420 234.570 33.920 234.830 ;
        LAYER Metal2 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  22.740 0.000 31.890 235.000 ;
        RECT  18.270 1.860 22.740 235.000 ;
        RECT  0.000 0.000 18.270 235.000 ;
        LAYER Via23 ;
        RECT  32.940 234.570 33.200 234.830 ;
        LAYER Metal3 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via34 ;
        RECT  32.420 234.570 33.920 234.830 ;
        LAYER Metal4 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via45 ;
        RECT  32.940 234.570 33.200 234.830 ;
        LAYER Metal5 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via56 ;
        RECT  32.370 234.520 33.970 234.880 ;
        LAYER Metal6 ;
        RECT  34.630 0.000 40.000 235.000 ;
        RECT  31.710 0.000 34.630 233.940 ;
        RECT  0.000 0.000 31.710 235.000 ;
    END
END PDIDGZ

MACRO PDO04CDG
    CLASS PAD ;
    FOREIGN PDO04CDG 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION OUTPUT ;
	AntennaDiffArea 2436.000000 ;
        PORT
        LAYER Metal1 ;
        RECT  18.550 0.000 22.460 1.580 ;
        LAYER Metal2 ;
        RECT  18.550 0.000 22.460 1.580 ;
        END
    END PAD
    PIN I
        DIRECTION INPUT ;
	AntennaGateArea 9.700000 ;
        PORT
        LAYER Metal1 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal2 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal3 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal4 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal5 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal6 ;
        RECT  32.170 234.400 34.170 235.000 ;
        END
    END I
    OBS
        LAYER Metal1 ;
        RECT  34.400 0.000 40.000 235.000 ;
        RECT  31.940 0.000 34.400 234.170 ;
        RECT  22.690 0.000 31.940 235.000 ;
        RECT  18.320 1.810 22.690 235.000 ;
        RECT  0.000 0.000 18.320 235.000 ;
        LAYER Via12 ;
        RECT  32.420 234.570 33.920 234.830 ;
        LAYER Metal2 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  22.740 0.000 31.890 235.000 ;
        RECT  18.270 1.860 22.740 235.000 ;
        RECT  0.000 0.000 18.270 235.000 ;
        LAYER Via23 ;
        RECT  32.940 234.570 33.200 234.830 ;
        LAYER Metal3 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via34 ;
        RECT  32.420 234.570 33.920 234.830 ;
        LAYER Metal4 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via45 ;
        RECT  32.940 234.570 33.200 234.830 ;
        LAYER Metal5 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  0.000 0.000 31.890 235.000 ;
        LAYER Via56 ;
        RECT  32.370 234.520 33.970 234.880 ;
        LAYER Metal6 ;
        RECT  34.630 0.000 40.000 235.000 ;
        RECT  31.710 0.000 34.630 233.940 ;
        RECT  0.000 0.000 31.710 235.000 ;
    END
END PDO04CDG

MACRO PFEED01
    CLASS PAD ;
    FOREIGN PFEED01 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.100 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 0.100 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 0.100 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 0.100 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 0.100 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 0.100 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 0.100 235.000 ;
    END
END PFEED01

MACRO PFEED1
    CLASS PAD ;
    FOREIGN PFEED1 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 1.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 1.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 1.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 1.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 1.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 1.000 235.000 ;
    END
END PFEED1

MACRO PFEED10
    CLASS PAD ;
    FOREIGN PFEED10 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 10.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 10.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 10.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 10.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 10.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 10.000 235.000 ;
    END
END PFEED10

MACRO PFEED2
    CLASS PAD ;
    FOREIGN PFEED2 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 2.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 2.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 2.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 2.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 2.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 2.000 235.000 ;
    END
END PFEED2

MACRO PFEED20
    CLASS PAD ;
    FOREIGN PFEED20 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 20.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 20.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 20.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 20.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 20.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 20.000 235.000 ;
    END
END PFEED20

MACRO PFEED35
    CLASS PAD ;
    FOREIGN PFEED35 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 35.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 35.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 35.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 35.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 35.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 35.000 235.000 ;
    END
END PFEED35

MACRO PFEED5
    CLASS PAD ;
    FOREIGN PFEED5 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 5.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 5.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 5.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 5.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 5.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 5.000 235.000 ;
    END
END PFEED5

MACRO PFEED50
    CLASS PAD ;
    FOREIGN PFEED50 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 50.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    OBS
        LAYER Metal1 ;
        RECT  0.000 0.000 50.000 235.000 ;
        LAYER Metal2 ;
        RECT  0.000 0.000 50.000 235.000 ;
        LAYER Metal3 ;
        RECT  0.000 0.000 50.000 235.000 ;
        LAYER Metal4 ;
        RECT  0.000 0.000 50.000 235.000 ;
        LAYER Metal5 ;
        RECT  0.000 0.000 50.000 235.000 ;
        LAYER Metal6 ;
        RECT  0.000 0.000 50.000 235.000 ;
    END
END PFEED50

MACRO PVDD1DGZ
    CLASS PAD POWER ;
    FOREIGN PVDD1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN VDD
        DIRECTION OUTPUT ;
	AntennaDiffArea 2616.960000 ;
        USE power ;
        PORT
	CLASS CORE ;
        LAYER Metal1 ;
        RECT  5.355 207.720 34.645 235.000 ;
        LAYER Metal2 ;
        RECT  5.355 207.720 34.645 235.000 ;
        LAYER Metal3 ;
        RECT  5.355 226.625 34.645 235.000 ;
        LAYER Metal4 ;
        RECT  5.355 226.625 34.645 235.000 ;
        LAYER Metal5 ;
        RECT  5.355 226.625 34.645 235.000 ;
        LAYER Metal6 ;
        RECT  5.355 226.625 34.645 235.000 ;
        END
    END VDD
    OBS
        LAYER Metal1 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 207.120 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via12 ;
        RECT  5.355 227.480 34.645 232.940 ;
        RECT  28.820 208.680 34.280 224.540 ;
        RECT  21.120 208.680 26.580 224.540 ;
        RECT  13.420 208.680 18.880 224.540 ;
        RECT  5.720 208.680 11.180 224.540 ;
        LAYER Metal2 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 207.120 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via23 ;
        RECT  34.170 234.570 34.485 234.830 ;
        RECT  6.165 226.960 34.170 234.830 ;
        RECT  5.830 226.960 6.165 233.460 ;
        LAYER Metal3 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 226.025 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via34 ;
        RECT  33.875 227.480 34.645 232.940 ;
        RECT  5.555 227.480 33.875 234.830 ;
        RECT  5.355 227.480 5.555 232.940 ;
        LAYER Metal4 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 226.025 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via45 ;
        RECT  34.170 234.570 34.485 234.830 ;
        RECT  6.165 226.960 34.170 234.830 ;
        RECT  5.830 226.960 6.165 233.460 ;
        LAYER Metal5 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 226.025 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via56 ;
        RECT  33.925 227.430 34.645 232.990 ;
        RECT  5.505 227.430 33.925 234.880 ;
        RECT  5.355 227.430 5.505 232.990 ;
        LAYER Metal6 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 226.025 ;
        RECT  0.000 0.000 4.755 235.000 ;
    END
END PVDD1DGZ

MACRO PVSS1DGZ
    CLASS PAD POWER ;
    FOREIGN PVSS1DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN VSS
        DIRECTION OUTPUT ;
	AntennaDiffArea 2616.960000 ;
        USE ground ;
        PORT
	CLASS CORE ;
        LAYER Metal1 ;
        RECT  5.355 207.720 34.645 235.000 ;
        LAYER Metal2 ;
        RECT  5.355 207.720 34.645 235.000 ;
        LAYER Metal3 ;
        RECT  5.355 234.400 34.645 235.000 ;
        LAYER Metal4 ;
        RECT  5.355 234.400 34.645 235.000 ;
        LAYER Metal5 ;
        RECT  5.355 234.400 34.645 235.000 ;
        LAYER Metal6 ;
        RECT  5.355 234.400 34.645 235.000 ;
        END
    END VSS
    OBS
        LAYER Metal1 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 207.120 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via12 ;
        RECT  28.820 208.680 34.280 224.540 ;
        RECT  6.350 227.480 33.650 232.940 ;
        RECT  21.120 208.680 26.580 224.540 ;
        RECT  13.420 208.680 18.880 224.540 ;
        RECT  5.720 208.680 11.180 224.540 ;
        LAYER Metal2 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 207.120 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via23 ;
        RECT  6.165 234.570 34.485 234.830 ;
        RECT  5.830 218.040 34.170 224.540 ;
        LAYER Metal3 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 233.800 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via34 ;
        RECT  5.555 234.570 33.875 234.830 ;
        LAYER Metal4 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 233.800 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via45 ;
        RECT  6.165 234.570 34.485 234.830 ;
        LAYER Metal5 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 233.800 ;
        RECT  0.000 0.000 4.755 235.000 ;
        LAYER Via56 ;
        RECT  5.505 234.520 33.925 234.880 ;
        LAYER Metal6 ;
        RECT  35.245 0.000 40.000 235.000 ;
        RECT  4.755 0.000 35.245 233.800 ;
        RECT  0.000 0.000 4.755 235.000 ;
    END
END PVSS1DGZ

MACRO PDB04DGZ
    CLASS PAD ;
    FOREIGN PDB04DGZ 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 40.000 BY 235.000 ;
    SYMMETRY x y r90 ;
    SITE pad ;
    PIN PAD
        DIRECTION INOUT ;
        PORT
        LAYER Metal1 ;
        RECT  18.550 0.000 22.460 1.580 ;
        LAYER Metal2 ;
        RECT  18.550 0.000 22.460 1.580 ;
        END
    END PAD
    PIN OEN
        DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  13.815 234.400 15.815 235.000 ;
        LAYER Metal2 ;
        RECT  13.815 234.400 15.815 235.000 ;
        LAYER Metal3 ;
        RECT  13.815 234.400 15.815 235.000 ;
        LAYER Metal4 ;
        RECT  13.815 234.400 15.815 235.000 ;
        LAYER Metal5 ;
        RECT  13.815 234.400 15.815 235.000 ;
        LAYER Metal6 ;
        RECT  13.815 234.400 15.815 235.000 ;
        END
    END OEN
    PIN I
        DIRECTION INPUT ;
        PORT
        LAYER Metal1 ;
        RECT  19.575 234.400 21.575 235.000 ;
        LAYER Metal2 ;
        RECT  19.575 234.400 21.575 235.000 ;
        LAYER Metal3 ;
        RECT  19.575 234.400 21.575 235.000 ;
        LAYER Metal4 ;
        RECT  19.575 234.400 21.575 235.000 ;
        LAYER Metal5 ;
        RECT  19.575 234.400 21.575 235.000 ;
        LAYER Metal6 ;
        RECT  19.575 234.400 21.575 235.000 ;
        END
    END I
    PIN C
        DIRECTION OUTPUT ;
        PORT
        LAYER Metal1 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal2 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal3 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal4 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal5 ;
        RECT  32.170 234.400 34.170 235.000 ;
        LAYER Metal6 ;
        RECT  32.170 234.400 34.170 235.000 ;
        END
    END C
    OBS
        LAYER Metal1 ;
        RECT  34.400 0.000 40.000 235.000 ;
        RECT  31.940 0.000 34.400 234.170 ;
        RECT  22.690 0.000 31.940 235.000 ;
        RECT  21.805 1.810 22.690 235.000 ;
        RECT  19.345 1.810 21.805 234.170 ;
        RECT  18.320 1.810 19.345 235.000 ;
        RECT  16.045 0.000 18.320 235.000 ;
        RECT  13.585 0.000 16.045 234.170 ;
        RECT  0.000 0.000 13.585 235.000 ;
        LAYER Via12 ;
        RECT  32.420 234.570 33.920 234.830 ;
        RECT  19.825 234.570 21.325 234.830 ;
        RECT  14.065 234.570 15.565 234.830 ;
        LAYER Metal2 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  22.740 0.000 31.890 235.000 ;
        RECT  21.855 1.860 22.740 235.000 ;
        RECT  19.295 1.860 21.855 234.120 ;
        RECT  18.270 1.860 19.295 235.000 ;
        RECT  16.095 0.000 18.270 235.000 ;
        RECT  13.535 0.000 16.095 234.120 ;
        RECT  0.000 0.000 13.535 235.000 ;
        LAYER Via23 ;
        RECT  32.940 234.570 33.200 234.830 ;
        RECT  20.345 234.570 20.605 234.830 ;
        RECT  14.585 234.570 14.845 234.830 ;
        LAYER Metal3 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  21.855 0.000 31.890 235.000 ;
        RECT  19.295 0.000 21.855 234.120 ;
        RECT  16.095 0.000 19.295 235.000 ;
        RECT  13.535 0.000 16.095 234.120 ;
        RECT  0.000 0.000 13.535 235.000 ;
        LAYER Via34 ;
        RECT  32.420 234.570 33.920 234.830 ;
        RECT  19.825 234.570 21.325 234.830 ;
        RECT  14.065 234.570 15.565 234.830 ;
        LAYER Metal4 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  21.855 0.000 31.890 235.000 ;
        RECT  19.295 0.000 21.855 234.120 ;
        RECT  16.095 0.000 19.295 235.000 ;
        RECT  13.535 0.000 16.095 234.120 ;
        RECT  0.000 0.000 13.535 235.000 ;
        LAYER Via45 ;
        RECT  32.940 234.570 33.200 234.830 ;
        RECT  20.345 234.570 20.605 234.830 ;
        RECT  14.585 234.570 14.845 234.830 ;
        LAYER Metal5 ;
        RECT  34.450 0.000 40.000 235.000 ;
        RECT  31.890 0.000 34.450 234.120 ;
        RECT  21.855 0.000 31.890 235.000 ;
        RECT  19.295 0.000 21.855 234.120 ;
        RECT  16.095 0.000 19.295 235.000 ;
        RECT  13.535 0.000 16.095 234.120 ;
        RECT  0.000 0.000 13.535 235.000 ;
        LAYER Via56 ;
        RECT  32.370 234.520 33.970 234.880 ;
        RECT  19.775 234.520 21.375 234.880 ;
        RECT  14.015 234.520 15.615 234.880 ;
        LAYER Metal6 ;
        RECT  34.630 0.000 40.000 235.000 ;
        RECT  31.710 0.000 34.630 233.940 ;
        RECT  22.035 0.000 31.710 235.000 ;
        RECT  19.115 0.000 22.035 233.940 ;
        RECT  16.275 0.000 19.115 235.000 ;
        RECT  13.355 0.000 16.275 233.940 ;
        RECT  0.000 0.000 13.355 235.000 ;
    END
END PDB04DGZ


MACRO ram_128x16A
  CLASS RING ;
  FOREIGN ram_128x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 593.82 BY 168.995 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 305.58 17.2 306.68 18.3 ;
      LAYER Metal2 ;
      RECT 305.58 17.2 306.68 18.3 ;
      LAYER Metal3 ;
      RECT 305.58 17.2 306.68 18.3 ;
      LAYER Metal4 ;
      RECT 305.58 17.2 306.68 18.3 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 301.92 17.2 303.02 18.3 ;
      LAYER Metal2 ;
      RECT 301.92 17.2 303.02 18.3 ;
      LAYER Metal3 ;
      RECT 301.92 17.2 303.02 18.3 ;
      LAYER Metal4 ;
      RECT 301.92 17.2 303.02 18.3 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 296.78 17.2 297.88 18.3 ;
      LAYER Metal2 ;
      RECT 296.78 17.2 297.88 18.3 ;
      LAYER Metal3 ;
      RECT 296.78 17.2 297.88 18.3 ;
      LAYER Metal4 ;
      RECT 296.78 17.2 297.88 18.3 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 293.12 17.2 294.22 18.3 ;
      LAYER Metal2 ;
      RECT 293.12 17.2 294.22 18.3 ;
      LAYER Metal3 ;
      RECT 293.12 17.2 294.22 18.3 ;
      LAYER Metal4 ;
      RECT 293.12 17.2 294.22 18.3 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 284.32 17.2 285.42 18.3 ;
      LAYER Metal2 ;
      RECT 284.32 17.2 285.42 18.3 ;
      LAYER Metal3 ;
      RECT 284.32 17.2 285.42 18.3 ;
      LAYER Metal4 ;
      RECT 284.32 17.2 285.42 18.3 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 279.18 17.2 280.28 18.3 ;
      LAYER Metal2 ;
      RECT 279.18 17.2 280.28 18.3 ;
      LAYER Metal3 ;
      RECT 279.18 17.2 280.28 18.3 ;
      LAYER Metal4 ;
      RECT 279.18 17.2 280.28 18.3 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 275.52 17.2 276.62 18.3 ;
      LAYER Metal2 ;
      RECT 275.52 17.2 276.62 18.3 ;
      LAYER Metal3 ;
      RECT 275.52 17.2 276.62 18.3 ;
      LAYER Metal4 ;
      RECT 275.52 17.2 276.62 18.3 ;
      END
    END A[6]
  PIN CEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 314.28 17.2 315.38 18.3 ;
      LAYER Metal2 ;
      RECT 314.28 17.2 315.38 18.3 ;
      LAYER Metal3 ;
      RECT 314.28 17.2 315.38 18.3 ;
      LAYER Metal4 ;
      RECT 314.28 17.2 315.38 18.3 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
      RECT 328.81 17.2 329.91 18.3 ;
      LAYER Metal2 ;
      RECT 328.81 17.2 329.91 18.3 ;
      LAYER Metal3 ;
      RECT 328.81 17.2 329.91 18.3 ;
      LAYER Metal4 ;
      RECT 328.81 17.2 329.91 18.3 ;
      END
    END CLK
  PIN D[0]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal2 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal3 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal4 ;
      RECT 45.46 17.2 46.56 18.3 ;
      END
    END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 415.08 17.2 416.18 18.3 ;
      LAYER Metal2 ;
      RECT 415.08 17.2 416.18 18.3 ;
      LAYER Metal3 ;
      RECT 415.08 17.2 416.18 18.3 ;
      LAYER Metal4 ;
      RECT 415.08 17.2 416.18 18.3 ;
      END
    END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 425.9 17.2 427 18.3 ;
      LAYER Metal2 ;
      RECT 425.9 17.2 427 18.3 ;
      LAYER Metal3 ;
      RECT 425.9 17.2 427 18.3 ;
      LAYER Metal4 ;
      RECT 425.9 17.2 427 18.3 ;
      END
    END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 475.76 17.2 476.86 18.3 ;
      LAYER Metal2 ;
      RECT 475.76 17.2 476.86 18.3 ;
      LAYER Metal3 ;
      RECT 475.76 17.2 476.86 18.3 ;
      LAYER Metal4 ;
      RECT 475.76 17.2 476.86 18.3 ;
      END
    END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 486.58 17.2 487.68 18.3 ;
      LAYER Metal2 ;
      RECT 486.58 17.2 487.68 18.3 ;
      LAYER Metal3 ;
      RECT 486.58 17.2 487.68 18.3 ;
      LAYER Metal4 ;
      RECT 486.58 17.2 487.68 18.3 ;
      END
    END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 536.44 17.2 537.54 18.3 ;
      LAYER Metal2 ;
      RECT 536.44 17.2 537.54 18.3 ;
      LAYER Metal3 ;
      RECT 536.44 17.2 537.54 18.3 ;
      LAYER Metal4 ;
      RECT 536.44 17.2 537.54 18.3 ;
      END
    END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 547.26 17.2 548.36 18.3 ;
      LAYER Metal2 ;
      RECT 547.26 17.2 548.36 18.3 ;
      LAYER Metal3 ;
      RECT 547.26 17.2 548.36 18.3 ;
      LAYER Metal4 ;
      RECT 547.26 17.2 548.36 18.3 ;
      END
    END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal2 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal3 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal4 ;
      RECT 56.28 17.2 57.38 18.3 ;
      END
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal2 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal3 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal4 ;
      RECT 106.14 17.2 107.24 18.3 ;
      END
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal2 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal3 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal4 ;
      RECT 116.96 17.2 118.06 18.3 ;
      END
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal2 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal3 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal4 ;
      RECT 166.82 17.2 167.92 18.3 ;
      END
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal2 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal3 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal4 ;
      RECT 177.64 17.2 178.74 18.3 ;
      END
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal2 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal3 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal4 ;
      RECT 227.5 17.2 228.6 18.3 ;
      END
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal2 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal3 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal4 ;
      RECT 238.32 17.2 239.42 18.3 ;
      END
    END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 354.4 17.2 355.5 18.3 ;
      LAYER Metal2 ;
      RECT 354.4 17.2 355.5 18.3 ;
      LAYER Metal3 ;
      RECT 354.4 17.2 355.5 18.3 ;
      LAYER Metal4 ;
      RECT 354.4 17.2 355.5 18.3 ;
      END
    END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 365.22 17.2 366.32 18.3 ;
      LAYER Metal2 ;
      RECT 365.22 17.2 366.32 18.3 ;
      LAYER Metal3 ;
      RECT 365.22 17.2 366.32 18.3 ;
      LAYER Metal4 ;
      RECT 365.22 17.2 366.32 18.3 ;
      END
    END D[9]
  PIN OEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 325.8 17.2 326.9 18.3 ;
      LAYER Metal2 ;
      RECT 325.8 17.2 326.9 18.3 ;
      LAYER Metal3 ;
      RECT 325.8 17.2 326.9 18.3 ;
      LAYER Metal4 ;
      RECT 325.8 17.2 326.9 18.3 ;
      END
    END OEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal2 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal3 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal4 ;
      RECT 39.98 17.2 41.08 18.3 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 409.8 17.2 410.9 18.3 ;
      LAYER Metal2 ;
      RECT 409.8 17.2 410.9 18.3 ;
      LAYER Metal3 ;
      RECT 409.8 17.2 410.9 18.3 ;
      LAYER Metal4 ;
      RECT 409.8 17.2 410.9 18.3 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 431.18 17.2 432.28 18.3 ;
      LAYER Metal2 ;
      RECT 431.18 17.2 432.28 18.3 ;
      LAYER Metal3 ;
      RECT 431.18 17.2 432.28 18.3 ;
      LAYER Metal4 ;
      RECT 431.18 17.2 432.28 18.3 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 470.48 17.2 471.58 18.3 ;
      LAYER Metal2 ;
      RECT 470.48 17.2 471.58 18.3 ;
      LAYER Metal3 ;
      RECT 470.48 17.2 471.58 18.3 ;
      LAYER Metal4 ;
      RECT 470.48 17.2 471.58 18.3 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 491.86 17.2 492.96 18.3 ;
      LAYER Metal2 ;
      RECT 491.86 17.2 492.96 18.3 ;
      LAYER Metal3 ;
      RECT 491.86 17.2 492.96 18.3 ;
      LAYER Metal4 ;
      RECT 491.86 17.2 492.96 18.3 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 531.16 17.2 532.26 18.3 ;
      LAYER Metal2 ;
      RECT 531.16 17.2 532.26 18.3 ;
      LAYER Metal3 ;
      RECT 531.16 17.2 532.26 18.3 ;
      LAYER Metal4 ;
      RECT 531.16 17.2 532.26 18.3 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 552.64 17.2 553.74 18.3 ;
      LAYER Metal2 ;
      RECT 552.64 17.2 553.74 18.3 ;
      LAYER Metal3 ;
      RECT 552.64 17.2 553.74 18.3 ;
      LAYER Metal4 ;
      RECT 552.64 17.2 553.74 18.3 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal2 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal3 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal4 ;
      RECT 61.56 17.2 62.66 18.3 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal2 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal3 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal4 ;
      RECT 100.86 17.2 101.96 18.3 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal2 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal3 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal4 ;
      RECT 122.24 17.2 123.34 18.3 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal2 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal3 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal4 ;
      RECT 161.54 17.2 162.64 18.3 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal2 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal3 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal4 ;
      RECT 182.92 17.2 184.02 18.3 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal2 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal3 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal4 ;
      RECT 222.22 17.2 223.32 18.3 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal2 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal3 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal4 ;
      RECT 243.6 17.2 244.7 18.3 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 349.12 17.2 350.22 18.3 ;
      LAYER Metal2 ;
      RECT 349.12 17.2 350.22 18.3 ;
      LAYER Metal3 ;
      RECT 349.12 17.2 350.22 18.3 ;
      LAYER Metal4 ;
      RECT 349.12 17.2 350.22 18.3 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 370.5 17.2 371.6 18.3 ;
      LAYER Metal2 ;
      RECT 370.5 17.2 371.6 18.3 ;
      LAYER Metal3 ;
      RECT 370.5 17.2 371.6 18.3 ;
      LAYER Metal4 ;
      RECT 370.5 17.2 371.6 18.3 ;
      END
    END Q[9]
  PIN WEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 317.16 17.2 318.26 18.3 ;
      LAYER Metal2 ;
      RECT 317.16 17.2 318.26 18.3 ;
      LAYER Metal3 ;
      RECT 317.16 17.2 318.26 18.3 ;
      LAYER Metal4 ;
      RECT 317.16 17.2 318.26 18.3 ;
      END
    END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 593.82 160.995 0 168.995 ;
      LAYER Metal5 ;
      RECT 0 0 593.82 8 ;
      LAYER Metal3 ;
      RECT 593.82 160.995 0 168.995 ;
      LAYER Metal3 ;
      RECT 0 0 593.82 8 ;
      LAYER Metal4 ;
      RECT 585.82 0 593.82 168.995 ;
      LAYER Metal4 ;
      RECT 0 168.995 8 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 585.22 152.395 8.6 160.395 ;
      LAYER Metal5 ;
      RECT 8.6 8.6 585.22 16.6 ;
      LAYER Metal3 ;
      RECT 585.22 152.395 8.6 160.395 ;
      LAYER Metal3 ;
      RECT 8.6 8.6 585.22 16.6 ;
      LAYER Metal4 ;
      RECT 577.22 8.6 585.22 160.395 ;
      LAYER Metal4 ;
      RECT 8.6 160.395 16.6 8.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Metal1 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Metal2 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Metal3 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Metal4 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Via12 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Via23 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Via34 ;
    RECT 17.2 17.2 576.62 151.795 ;
    LAYER Via34 ;
    RECT 577.45 152.625 584.99 160.165 ;
    LAYER Via34 ;
    RECT 8.83 8.83 16.37 16.37 ;
    LAYER Via34 ;
    RECT 577.45 8.83 584.99 16.37 ;
    LAYER Via34 ;
    RECT 8.83 152.625 16.37 160.165 ;
    LAYER Via34 ;
    RECT 586.05 161.225 593.59 168.765 ;
    LAYER Via34 ;
    RECT 0.23 0.23 7.77 7.77 ;
    LAYER Via34 ;
    RECT 586.05 0.23 593.59 7.77 ;
    LAYER Via34 ;
    RECT 0.23 161.225 7.77 168.765 ;
    LAYER Metal4 ;
    RECT 18.62 151.795 19.7 168.995 ;
    LAYER Metal4 ;
    RECT 24.1 151.795 25.26 168.995 ;
    LAYER Metal4 ;
    RECT 26.06 151.795 27.22 168.995 ;
    LAYER Metal4 ;
    RECT 31.46 151.795 32.62 168.995 ;
    LAYER Metal4 ;
    RECT 33.42 151.795 34.58 168.995 ;
    LAYER Metal4 ;
    RECT 38.82 151.795 39.98 168.995 ;
    LAYER Metal4 ;
    RECT 40.78 151.795 41.94 168.995 ;
    LAYER Metal4 ;
    RECT 46.18 151.795 47.34 168.995 ;
    LAYER Metal4 ;
    RECT 48.14 151.795 49.3 168.995 ;
    LAYER Metal4 ;
    RECT 53.54 151.795 54.7 168.995 ;
    LAYER Metal4 ;
    RECT 55.5 151.795 56.66 168.995 ;
    LAYER Metal4 ;
    RECT 60.9 151.795 62.06 168.995 ;
    LAYER Metal4 ;
    RECT 62.86 151.795 64.02 168.995 ;
    LAYER Metal4 ;
    RECT 68.26 151.795 69.42 168.995 ;
    LAYER Metal4 ;
    RECT 70.22 151.795 71.38 168.995 ;
    LAYER Metal4 ;
    RECT 75.62 151.795 76.78 168.995 ;
    LAYER Metal4 ;
    RECT 77.58 151.795 78.74 168.995 ;
    LAYER Metal4 ;
    RECT 84.78 151.795 85.94 168.995 ;
    LAYER Metal4 ;
    RECT 86.74 151.795 87.9 168.995 ;
    LAYER Metal4 ;
    RECT 92.14 151.795 93.3 168.995 ;
    LAYER Metal4 ;
    RECT 94.1 151.795 95.26 168.995 ;
    LAYER Metal4 ;
    RECT 99.5 151.795 100.66 168.995 ;
    LAYER Metal4 ;
    RECT 101.46 151.795 102.62 168.995 ;
    LAYER Metal4 ;
    RECT 106.86 151.795 108.02 168.995 ;
    LAYER Metal4 ;
    RECT 108.82 151.795 109.98 168.995 ;
    LAYER Metal4 ;
    RECT 114.22 151.795 115.38 168.995 ;
    LAYER Metal4 ;
    RECT 116.18 151.795 117.34 168.995 ;
    LAYER Metal4 ;
    RECT 121.58 151.795 122.74 168.995 ;
    LAYER Metal4 ;
    RECT 123.54 151.795 124.7 168.995 ;
    LAYER Metal4 ;
    RECT 128.94 151.795 130.1 168.995 ;
    LAYER Metal4 ;
    RECT 130.9 151.795 132.06 168.995 ;
    LAYER Metal4 ;
    RECT 136.3 151.795 137.46 168.995 ;
    LAYER Metal4 ;
    RECT 138.26 151.795 139.42 168.995 ;
    LAYER Metal4 ;
    RECT 145.46 151.795 146.62 168.995 ;
    LAYER Metal4 ;
    RECT 147.42 151.795 148.58 168.995 ;
    LAYER Metal4 ;
    RECT 152.82 151.795 153.98 168.995 ;
    LAYER Metal4 ;
    RECT 154.78 151.795 155.94 168.995 ;
    LAYER Metal4 ;
    RECT 160.18 151.795 161.34 168.995 ;
    LAYER Metal4 ;
    RECT 162.14 151.795 163.3 168.995 ;
    LAYER Metal4 ;
    RECT 167.54 151.795 168.7 168.995 ;
    LAYER Metal4 ;
    RECT 169.5 151.795 170.66 168.995 ;
    LAYER Metal4 ;
    RECT 174.9 151.795 176.06 168.995 ;
    LAYER Metal4 ;
    RECT 176.86 151.795 178.02 168.995 ;
    LAYER Metal4 ;
    RECT 182.26 151.795 183.42 168.995 ;
    LAYER Metal4 ;
    RECT 184.22 151.795 185.38 168.995 ;
    LAYER Metal4 ;
    RECT 189.62 151.795 190.78 168.995 ;
    LAYER Metal4 ;
    RECT 191.58 151.795 192.74 168.995 ;
    LAYER Metal4 ;
    RECT 196.98 151.795 198.14 168.995 ;
    LAYER Metal4 ;
    RECT 198.94 151.795 200.1 168.995 ;
    LAYER Metal4 ;
    RECT 206.14 151.795 207.3 168.995 ;
    LAYER Metal4 ;
    RECT 208.1 151.795 209.26 168.995 ;
    LAYER Metal4 ;
    RECT 213.5 151.795 214.66 168.995 ;
    LAYER Metal4 ;
    RECT 215.46 151.795 216.62 168.995 ;
    LAYER Metal4 ;
    RECT 220.86 151.795 222.02 168.995 ;
    LAYER Metal4 ;
    RECT 222.82 151.795 223.98 168.995 ;
    LAYER Metal4 ;
    RECT 228.22 151.795 229.38 168.995 ;
    LAYER Metal4 ;
    RECT 230.18 151.795 231.34 168.995 ;
    LAYER Metal4 ;
    RECT 235.58 151.795 236.74 168.995 ;
    LAYER Metal4 ;
    RECT 237.54 151.795 238.7 168.995 ;
    LAYER Metal4 ;
    RECT 242.94 151.795 244.1 168.995 ;
    LAYER Metal4 ;
    RECT 244.9 151.795 246.06 168.995 ;
    LAYER Metal4 ;
    RECT 250.3 151.795 251.46 168.995 ;
    LAYER Metal4 ;
    RECT 252.26 151.795 253.42 168.995 ;
    LAYER Metal4 ;
    RECT 257.66 151.795 258.82 168.995 ;
    LAYER Metal4 ;
    RECT 259.62 151.795 260.78 168.995 ;
    LAYER Metal4 ;
    RECT 264.96 151.795 266.64 168.995 ;
    LAYER Metal4 ;
    RECT 269.36 151.795 271.04 168.995 ;
    LAYER Metal4 ;
    RECT 273.76 151.795 275.44 168.995 ;
    LAYER Metal4 ;
    RECT 278.16 151.795 279.84 168.995 ;
    LAYER Metal4 ;
    RECT 282.56 151.795 284.24 168.995 ;
    LAYER Metal4 ;
    RECT 286.96 151.795 288.64 168.995 ;
    LAYER Metal4 ;
    RECT 291.36 151.795 293.04 168.995 ;
    LAYER Metal4 ;
    RECT 295.76 151.795 297.44 168.995 ;
    LAYER Metal4 ;
    RECT 300.16 151.795 301.84 168.995 ;
    LAYER Metal4 ;
    RECT 304.56 151.795 306.24 168.995 ;
    LAYER Metal4 ;
    RECT 310.32 151.795 311.52 168.995 ;
    LAYER Metal4 ;
    RECT 315.26 151.795 317.28 168.995 ;
    LAYER Metal4 ;
    RECT 321.02 151.795 323.04 168.995 ;
    LAYER Metal4 ;
    RECT 325.72 151.795 327 168.995 ;
    LAYER Metal4 ;
    RECT 329.3 151.795 330.74 168.995 ;
    LAYER Metal4 ;
    RECT 333.04 151.795 334.2 168.995 ;
    LAYER Metal4 ;
    RECT 335 151.795 336.16 168.995 ;
    LAYER Metal4 ;
    RECT 340.4 151.795 341.56 168.995 ;
    LAYER Metal4 ;
    RECT 342.36 151.795 343.52 168.995 ;
    LAYER Metal4 ;
    RECT 347.76 151.795 348.92 168.995 ;
    LAYER Metal4 ;
    RECT 349.72 151.795 350.88 168.995 ;
    LAYER Metal4 ;
    RECT 355.12 151.795 356.28 168.995 ;
    LAYER Metal4 ;
    RECT 357.08 151.795 358.24 168.995 ;
    LAYER Metal4 ;
    RECT 362.48 151.795 363.64 168.995 ;
    LAYER Metal4 ;
    RECT 364.44 151.795 365.6 168.995 ;
    LAYER Metal4 ;
    RECT 369.84 151.795 371 168.995 ;
    LAYER Metal4 ;
    RECT 371.8 151.795 372.96 168.995 ;
    LAYER Metal4 ;
    RECT 377.2 151.795 378.36 168.995 ;
    LAYER Metal4 ;
    RECT 379.16 151.795 380.32 168.995 ;
    LAYER Metal4 ;
    RECT 384.56 151.795 385.72 168.995 ;
    LAYER Metal4 ;
    RECT 386.52 151.795 387.68 168.995 ;
    LAYER Metal4 ;
    RECT 393.72 151.795 394.88 168.995 ;
    LAYER Metal4 ;
    RECT 395.68 151.795 396.84 168.995 ;
    LAYER Metal4 ;
    RECT 401.08 151.795 402.24 168.995 ;
    LAYER Metal4 ;
    RECT 403.04 151.795 404.2 168.995 ;
    LAYER Metal4 ;
    RECT 408.44 151.795 409.6 168.995 ;
    LAYER Metal4 ;
    RECT 410.4 151.795 411.56 168.995 ;
    LAYER Metal4 ;
    RECT 415.8 151.795 416.96 168.995 ;
    LAYER Metal4 ;
    RECT 417.76 151.795 418.92 168.995 ;
    LAYER Metal4 ;
    RECT 423.16 151.795 424.32 168.995 ;
    LAYER Metal4 ;
    RECT 425.12 151.795 426.28 168.995 ;
    LAYER Metal4 ;
    RECT 430.52 151.795 431.68 168.995 ;
    LAYER Metal4 ;
    RECT 432.48 151.795 433.64 168.995 ;
    LAYER Metal4 ;
    RECT 437.88 151.795 439.04 168.995 ;
    LAYER Metal4 ;
    RECT 439.84 151.795 441 168.995 ;
    LAYER Metal4 ;
    RECT 445.24 151.795 446.4 168.995 ;
    LAYER Metal4 ;
    RECT 447.2 151.795 448.36 168.995 ;
    LAYER Metal4 ;
    RECT 454.4 151.795 455.56 168.995 ;
    LAYER Metal4 ;
    RECT 456.36 151.795 457.52 168.995 ;
    LAYER Metal4 ;
    RECT 461.76 151.795 462.92 168.995 ;
    LAYER Metal4 ;
    RECT 463.72 151.795 464.88 168.995 ;
    LAYER Metal4 ;
    RECT 469.12 151.795 470.28 168.995 ;
    LAYER Metal4 ;
    RECT 471.08 151.795 472.24 168.995 ;
    LAYER Metal4 ;
    RECT 476.48 151.795 477.64 168.995 ;
    LAYER Metal4 ;
    RECT 478.44 151.795 479.6 168.995 ;
    LAYER Metal4 ;
    RECT 483.84 151.795 485 168.995 ;
    LAYER Metal4 ;
    RECT 485.8 151.795 486.96 168.995 ;
    LAYER Metal4 ;
    RECT 491.2 151.795 492.36 168.995 ;
    LAYER Metal4 ;
    RECT 493.16 151.795 494.32 168.995 ;
    LAYER Metal4 ;
    RECT 498.56 151.795 499.72 168.995 ;
    LAYER Metal4 ;
    RECT 500.52 151.795 501.68 168.995 ;
    LAYER Metal4 ;
    RECT 505.92 151.795 507.08 168.995 ;
    LAYER Metal4 ;
    RECT 507.88 151.795 509.04 168.995 ;
    LAYER Metal4 ;
    RECT 515.08 151.795 516.24 168.995 ;
    LAYER Metal4 ;
    RECT 517.04 151.795 518.2 168.995 ;
    LAYER Metal4 ;
    RECT 522.44 151.795 523.6 168.995 ;
    LAYER Metal4 ;
    RECT 524.4 151.795 525.56 168.995 ;
    LAYER Metal4 ;
    RECT 529.8 151.795 530.96 168.995 ;
    LAYER Metal4 ;
    RECT 531.76 151.795 532.92 168.995 ;
    LAYER Metal4 ;
    RECT 537.16 151.795 538.32 168.995 ;
    LAYER Metal4 ;
    RECT 539.12 151.795 540.28 168.995 ;
    LAYER Metal4 ;
    RECT 544.52 151.795 545.68 168.995 ;
    LAYER Metal4 ;
    RECT 546.48 151.795 547.64 168.995 ;
    LAYER Metal4 ;
    RECT 551.88 151.795 553.04 168.995 ;
    LAYER Metal4 ;
    RECT 553.84 151.795 555 168.995 ;
    LAYER Metal4 ;
    RECT 559.24 151.795 560.4 168.995 ;
    LAYER Metal4 ;
    RECT 561.2 151.795 562.36 168.995 ;
    LAYER Metal4 ;
    RECT 566.6 151.795 567.76 168.995 ;
    LAYER Metal4 ;
    RECT 568.56 151.795 569.72 168.995 ;
    LAYER Metal4 ;
    RECT 574.12 151.795 575.2 168.995 ;
    LAYER Metal4 ;
    RECT 18.02 17.2 19.12 0 ;
    LAYER Metal4 ;
    RECT 24.1 17.2 27.22 0 ;
    LAYER Metal4 ;
    RECT 31.46 17.2 34.58 0 ;
    LAYER Metal4 ;
    RECT 38.18 17.2 39.52 0 ;
    LAYER Metal4 ;
    RECT 47.02 17.2 49.4 0 ;
    LAYER Metal4 ;
    RECT 53.44 17.2 55.82 0 ;
    LAYER Metal4 ;
    RECT 63.32 17.2 64.66 0 ;
    LAYER Metal4 ;
    RECT 68.26 17.2 71.38 0 ;
    LAYER Metal4 ;
    RECT 75.62 17.2 78.74 0 ;
    LAYER Metal4 ;
    RECT 84.78 17.2 87.9 0 ;
    LAYER Metal4 ;
    RECT 92.14 17.2 95.26 0 ;
    LAYER Metal4 ;
    RECT 98.86 17.2 100.2 0 ;
    LAYER Metal4 ;
    RECT 107.7 17.2 110.08 0 ;
    LAYER Metal4 ;
    RECT 114.12 17.2 116.5 0 ;
    LAYER Metal4 ;
    RECT 124 17.2 125.34 0 ;
    LAYER Metal4 ;
    RECT 128.94 17.2 132.06 0 ;
    LAYER Metal4 ;
    RECT 136.3 17.2 139.42 0 ;
    LAYER Metal4 ;
    RECT 145.46 17.2 148.58 0 ;
    LAYER Metal4 ;
    RECT 152.82 17.2 155.94 0 ;
    LAYER Metal4 ;
    RECT 159.54 17.2 160.88 0 ;
    LAYER Metal4 ;
    RECT 168.38 17.2 170.76 0 ;
    LAYER Metal4 ;
    RECT 174.8 17.2 177.18 0 ;
    LAYER Metal4 ;
    RECT 184.68 17.2 186.02 0 ;
    LAYER Metal4 ;
    RECT 189.62 17.2 192.74 0 ;
    LAYER Metal4 ;
    RECT 196.98 17.2 200.1 0 ;
    LAYER Metal4 ;
    RECT 206.14 17.2 209.26 0 ;
    LAYER Metal4 ;
    RECT 213.5 17.2 216.62 0 ;
    LAYER Metal4 ;
    RECT 220.22 17.2 221.56 0 ;
    LAYER Metal4 ;
    RECT 229.06 17.2 231.44 0 ;
    LAYER Metal4 ;
    RECT 235.48 17.2 237.86 0 ;
    LAYER Metal4 ;
    RECT 245.36 17.2 246.7 0 ;
    LAYER Metal4 ;
    RECT 250.3 17.2 253.42 0 ;
    LAYER Metal4 ;
    RECT 257.66 17.2 260.78 0 ;
    LAYER Metal4 ;
    RECT 270.58 17.2 274.38 0 ;
    LAYER Metal4 ;
    RECT 281.48 17.2 283.12 0 ;
    LAYER Metal4 ;
    RECT 288.18 17.2 291.98 0 ;
    LAYER Metal4 ;
    RECT 299.08 17.2 300.72 0 ;
    LAYER Metal4 ;
    RECT 308.43 17.2 308.97 0 ;
    LAYER Metal4 ;
    RECT 310.01 17.2 311.01 0 ;
    LAYER Metal4 ;
    RECT 315.84 17.2 316.7 0 ;
    LAYER Metal4 ;
    RECT 321.6 17.2 322.46 0 ;
    LAYER Metal4 ;
    RECT 333.04 17.2 336.16 0 ;
    LAYER Metal4 ;
    RECT 340.4 17.2 343.52 0 ;
    LAYER Metal4 ;
    RECT 347.12 17.2 348.46 0 ;
    LAYER Metal4 ;
    RECT 355.96 17.2 358.34 0 ;
    LAYER Metal4 ;
    RECT 362.38 17.2 364.76 0 ;
    LAYER Metal4 ;
    RECT 372.26 17.2 373.6 0 ;
    LAYER Metal4 ;
    RECT 377.2 17.2 380.32 0 ;
    LAYER Metal4 ;
    RECT 384.56 17.2 387.68 0 ;
    LAYER Metal4 ;
    RECT 393.72 17.2 396.84 0 ;
    LAYER Metal4 ;
    RECT 401.08 17.2 404.2 0 ;
    LAYER Metal4 ;
    RECT 407.8 17.2 409.14 0 ;
    LAYER Metal4 ;
    RECT 416.64 17.2 419.02 0 ;
    LAYER Metal4 ;
    RECT 423.06 17.2 425.44 0 ;
    LAYER Metal4 ;
    RECT 432.94 17.2 434.28 0 ;
    LAYER Metal4 ;
    RECT 437.88 17.2 441 0 ;
    LAYER Metal4 ;
    RECT 445.24 17.2 448.36 0 ;
    LAYER Metal4 ;
    RECT 454.4 17.2 457.52 0 ;
    LAYER Metal4 ;
    RECT 461.76 17.2 464.88 0 ;
    LAYER Metal4 ;
    RECT 468.48 17.2 469.82 0 ;
    LAYER Metal4 ;
    RECT 477.32 17.2 479.7 0 ;
    LAYER Metal4 ;
    RECT 483.74 17.2 486.12 0 ;
    LAYER Metal4 ;
    RECT 493.62 17.2 494.96 0 ;
    LAYER Metal4 ;
    RECT 498.56 17.2 501.68 0 ;
    LAYER Metal4 ;
    RECT 505.92 17.2 509.04 0 ;
    LAYER Metal4 ;
    RECT 515.08 17.2 518.2 0 ;
    LAYER Metal4 ;
    RECT 522.44 17.2 525.56 0 ;
    LAYER Metal4 ;
    RECT 529.16 17.2 530.5 0 ;
    LAYER Metal4 ;
    RECT 538 17.2 540.38 0 ;
    LAYER Metal4 ;
    RECT 544.42 17.2 546.8 0 ;
    LAYER Metal4 ;
    RECT 554.3 17.2 555.64 0 ;
    LAYER Metal4 ;
    RECT 559.24 17.2 562.36 0 ;
    LAYER Metal4 ;
    RECT 566.6 17.2 569.72 0 ;
    LAYER Metal4 ;
    RECT 574.7 17.2 575.8 0 ;
    LAYER Metal3 ;
    RECT 576.62 22.22 593.82 23.22 ;
    LAYER Metal3 ;
    RECT 576.62 35.14 593.82 36.04 ;
    LAYER Metal3 ;
    RECT 576.62 48.245 593.82 48.845 ;
    LAYER Metal3 ;
    RECT 576.62 52.605 593.82 53.505 ;
    LAYER Metal3 ;
    RECT 576.62 73.205 593.82 73.805 ;
    LAYER Metal3 ;
    RECT 576.62 82.685 593.82 84.285 ;
    LAYER Metal3 ;
    RECT 576.62 90.11 593.82 94.61 ;
    LAYER Metal3 ;
    RECT 576.62 95.21 593.82 103.61 ;
    LAYER Metal3 ;
    RECT 576.62 105.875 593.82 109.575 ;
    LAYER Metal3 ;
    RECT 576.62 110.19 593.82 114.19 ;
    LAYER Metal3 ;
    RECT 576.62 123.595 593.82 124.495 ;
    LAYER Metal3 ;
    RECT 576.62 128.655 593.82 129.555 ;
    LAYER Metal3 ;
    RECT 576.62 133.715 593.82 134.615 ;
    LAYER Metal3 ;
    RECT 576.62 138.775 593.82 139.675 ;
    LAYER Metal3 ;
    RECT 576.62 144.105 593.82 145.005 ;
    LAYER Metal3 ;
    RECT 576.62 148.005 593.82 148.905 ;
    LAYER Metal3 ;
    RECT 17.2 22.22 0 23.22 ;
    LAYER Metal3 ;
    RECT 17.2 35.14 0 36.04 ;
    LAYER Metal3 ;
    RECT 17.2 48.245 0 48.845 ;
    LAYER Metal3 ;
    RECT 17.2 52.605 0 53.505 ;
    LAYER Metal3 ;
    RECT 17.2 73.205 0 73.805 ;
    LAYER Metal3 ;
    RECT 17.2 82.685 0 84.285 ;
    LAYER Metal3 ;
    RECT 17.2 90.11 0 94.61 ;
    LAYER Metal3 ;
    RECT 17.2 95.21 0 103.61 ;
    LAYER Metal3 ;
    RECT 17.2 105.875 0 109.575 ;
    LAYER Metal3 ;
    RECT 17.2 110.19 0 114.19 ;
    LAYER Metal3 ;
    RECT 17.2 123.595 0 124.495 ;
    LAYER Metal3 ;
    RECT 17.2 128.655 0 129.555 ;
    LAYER Metal3 ;
    RECT 17.2 133.715 0 134.615 ;
    LAYER Metal3 ;
    RECT 17.2 138.775 0 139.675 ;
    LAYER Metal3 ;
    RECT 17.2 144.105 0 145.005 ;
    LAYER Metal3 ;
    RECT 17.2 148.005 0 148.905 ;
    LAYER Metal4 ;
    RECT 20.42 151.795 21.7 160.395 ;
    LAYER Metal4 ;
    RECT 22.38 151.795 23.54 160.395 ;
    LAYER Metal4 ;
    RECT 27.78 151.795 28.94 160.395 ;
    LAYER Metal4 ;
    RECT 29.74 151.795 30.9 160.395 ;
    LAYER Metal4 ;
    RECT 35.14 151.795 36.3 160.395 ;
    LAYER Metal4 ;
    RECT 37.1 151.795 38.26 160.395 ;
    LAYER Metal4 ;
    RECT 42.5 151.795 43.66 160.395 ;
    LAYER Metal4 ;
    RECT 44.46 151.795 45.62 160.395 ;
    LAYER Metal4 ;
    RECT 49.86 151.795 51.02 160.395 ;
    LAYER Metal4 ;
    RECT 51.82 151.795 52.98 160.395 ;
    LAYER Metal4 ;
    RECT 57.22 151.795 58.38 160.395 ;
    LAYER Metal4 ;
    RECT 59.18 151.795 60.34 160.395 ;
    LAYER Metal4 ;
    RECT 64.58 151.795 65.74 160.395 ;
    LAYER Metal4 ;
    RECT 66.54 151.795 67.7 160.395 ;
    LAYER Metal4 ;
    RECT 71.94 151.795 73.1 160.395 ;
    LAYER Metal4 ;
    RECT 73.9 151.795 75.06 160.395 ;
    LAYER Metal4 ;
    RECT 79.3 151.795 80.46 160.395 ;
    LAYER Metal4 ;
    RECT 81.21 151.795 82.31 160.395 ;
    LAYER Metal4 ;
    RECT 83.06 151.795 84.22 160.395 ;
    LAYER Metal4 ;
    RECT 88.46 151.795 89.62 160.395 ;
    LAYER Metal4 ;
    RECT 90.42 151.795 91.58 160.395 ;
    LAYER Metal4 ;
    RECT 95.82 151.795 96.98 160.395 ;
    LAYER Metal4 ;
    RECT 97.78 151.795 98.94 160.395 ;
    LAYER Metal4 ;
    RECT 103.18 151.795 104.34 160.395 ;
    LAYER Metal4 ;
    RECT 105.14 151.795 106.3 160.395 ;
    LAYER Metal4 ;
    RECT 110.54 151.795 111.7 160.395 ;
    LAYER Metal4 ;
    RECT 112.5 151.795 113.66 160.395 ;
    LAYER Metal4 ;
    RECT 117.9 151.795 119.06 160.395 ;
    LAYER Metal4 ;
    RECT 119.86 151.795 121.02 160.395 ;
    LAYER Metal4 ;
    RECT 125.26 151.795 126.42 160.395 ;
    LAYER Metal4 ;
    RECT 127.22 151.795 128.38 160.395 ;
    LAYER Metal4 ;
    RECT 132.62 151.795 133.78 160.395 ;
    LAYER Metal4 ;
    RECT 134.58 151.795 135.74 160.395 ;
    LAYER Metal4 ;
    RECT 139.98 151.795 141.14 160.395 ;
    LAYER Metal4 ;
    RECT 141.89 151.795 142.99 160.395 ;
    LAYER Metal4 ;
    RECT 143.74 151.795 144.9 160.395 ;
    LAYER Metal4 ;
    RECT 149.14 151.795 150.3 160.395 ;
    LAYER Metal4 ;
    RECT 151.1 151.795 152.26 160.395 ;
    LAYER Metal4 ;
    RECT 156.5 151.795 157.66 160.395 ;
    LAYER Metal4 ;
    RECT 158.46 151.795 159.62 160.395 ;
    LAYER Metal4 ;
    RECT 163.86 151.795 165.02 160.395 ;
    LAYER Metal4 ;
    RECT 165.82 151.795 166.98 160.395 ;
    LAYER Metal4 ;
    RECT 171.22 151.795 172.38 160.395 ;
    LAYER Metal4 ;
    RECT 173.18 151.795 174.34 160.395 ;
    LAYER Metal4 ;
    RECT 178.58 151.795 179.74 160.395 ;
    LAYER Metal4 ;
    RECT 180.54 151.795 181.7 160.395 ;
    LAYER Metal4 ;
    RECT 185.94 151.795 187.1 160.395 ;
    LAYER Metal4 ;
    RECT 187.9 151.795 189.06 160.395 ;
    LAYER Metal4 ;
    RECT 193.3 151.795 194.46 160.395 ;
    LAYER Metal4 ;
    RECT 195.26 151.795 196.42 160.395 ;
    LAYER Metal4 ;
    RECT 200.66 151.795 201.82 160.395 ;
    LAYER Metal4 ;
    RECT 202.57 151.795 203.67 160.395 ;
    LAYER Metal4 ;
    RECT 204.42 151.795 205.58 160.395 ;
    LAYER Metal4 ;
    RECT 209.82 151.795 210.98 160.395 ;
    LAYER Metal4 ;
    RECT 211.78 151.795 212.94 160.395 ;
    LAYER Metal4 ;
    RECT 217.18 151.795 218.34 160.395 ;
    LAYER Metal4 ;
    RECT 219.14 151.795 220.3 160.395 ;
    LAYER Metal4 ;
    RECT 224.54 151.795 225.7 160.395 ;
    LAYER Metal4 ;
    RECT 226.5 151.795 227.66 160.395 ;
    LAYER Metal4 ;
    RECT 231.9 151.795 233.06 160.395 ;
    LAYER Metal4 ;
    RECT 233.86 151.795 235.02 160.395 ;
    LAYER Metal4 ;
    RECT 239.26 151.795 240.42 160.395 ;
    LAYER Metal4 ;
    RECT 241.22 151.795 242.38 160.395 ;
    LAYER Metal4 ;
    RECT 246.62 151.795 247.78 160.395 ;
    LAYER Metal4 ;
    RECT 248.58 151.795 249.74 160.395 ;
    LAYER Metal4 ;
    RECT 253.98 151.795 255.14 160.395 ;
    LAYER Metal4 ;
    RECT 255.94 151.795 257.1 160.395 ;
    LAYER Metal4 ;
    RECT 261.34 151.795 262.5 160.395 ;
    LAYER Metal4 ;
    RECT 263.25 151.795 264.35 160.395 ;
    LAYER Metal4 ;
    RECT 267.1 151.795 268.9 160.395 ;
    LAYER Metal4 ;
    RECT 271.56 151.795 273.24 160.395 ;
    LAYER Metal4 ;
    RECT 275.96 151.795 277.64 160.395 ;
    LAYER Metal4 ;
    RECT 280.36 151.795 282.04 160.395 ;
    LAYER Metal4 ;
    RECT 284.76 151.795 286.44 160.395 ;
    LAYER Metal4 ;
    RECT 289.16 151.795 290.84 160.395 ;
    LAYER Metal4 ;
    RECT 293.56 151.795 295.24 160.395 ;
    LAYER Metal4 ;
    RECT 297.96 151.795 299.64 160.395 ;
    LAYER Metal4 ;
    RECT 302.36 151.795 304.04 160.395 ;
    LAYER Metal4 ;
    RECT 306.7 151.795 309.7 160.395 ;
    LAYER Metal4 ;
    RECT 312.38 151.795 314.4 160.395 ;
    LAYER Metal4 ;
    RECT 318.14 151.795 320.16 160.395 ;
    LAYER Metal4 ;
    RECT 323.9 151.795 325.1 160.395 ;
    LAYER Metal4 ;
    RECT 327.56 151.795 328.84 160.395 ;
    LAYER Metal4 ;
    RECT 331.32 151.795 332.48 160.395 ;
    LAYER Metal4 ;
    RECT 336.72 151.795 337.88 160.395 ;
    LAYER Metal4 ;
    RECT 338.68 151.795 339.84 160.395 ;
    LAYER Metal4 ;
    RECT 344.08 151.795 345.24 160.395 ;
    LAYER Metal4 ;
    RECT 346.04 151.795 347.2 160.395 ;
    LAYER Metal4 ;
    RECT 351.44 151.795 352.6 160.395 ;
    LAYER Metal4 ;
    RECT 353.4 151.795 354.56 160.395 ;
    LAYER Metal4 ;
    RECT 358.8 151.795 359.96 160.395 ;
    LAYER Metal4 ;
    RECT 360.76 151.795 361.92 160.395 ;
    LAYER Metal4 ;
    RECT 366.16 151.795 367.32 160.395 ;
    LAYER Metal4 ;
    RECT 368.12 151.795 369.28 160.395 ;
    LAYER Metal4 ;
    RECT 373.52 151.795 374.68 160.395 ;
    LAYER Metal4 ;
    RECT 375.48 151.795 376.64 160.395 ;
    LAYER Metal4 ;
    RECT 380.88 151.795 382.04 160.395 ;
    LAYER Metal4 ;
    RECT 382.84 151.795 384 160.395 ;
    LAYER Metal4 ;
    RECT 388.24 151.795 389.4 160.395 ;
    LAYER Metal4 ;
    RECT 390.15 151.795 391.25 160.395 ;
    LAYER Metal4 ;
    RECT 392 151.795 393.16 160.395 ;
    LAYER Metal4 ;
    RECT 397.4 151.795 398.56 160.395 ;
    LAYER Metal4 ;
    RECT 399.36 151.795 400.52 160.395 ;
    LAYER Metal4 ;
    RECT 404.76 151.795 405.92 160.395 ;
    LAYER Metal4 ;
    RECT 406.72 151.795 407.88 160.395 ;
    LAYER Metal4 ;
    RECT 412.12 151.795 413.28 160.395 ;
    LAYER Metal4 ;
    RECT 414.08 151.795 415.24 160.395 ;
    LAYER Metal4 ;
    RECT 419.48 151.795 420.64 160.395 ;
    LAYER Metal4 ;
    RECT 421.44 151.795 422.6 160.395 ;
    LAYER Metal4 ;
    RECT 426.84 151.795 428 160.395 ;
    LAYER Metal4 ;
    RECT 428.8 151.795 429.96 160.395 ;
    LAYER Metal4 ;
    RECT 434.2 151.795 435.36 160.395 ;
    LAYER Metal4 ;
    RECT 436.16 151.795 437.32 160.395 ;
    LAYER Metal4 ;
    RECT 441.56 151.795 442.72 160.395 ;
    LAYER Metal4 ;
    RECT 443.52 151.795 444.68 160.395 ;
    LAYER Metal4 ;
    RECT 448.92 151.795 450.08 160.395 ;
    LAYER Metal4 ;
    RECT 450.83 151.795 451.93 160.395 ;
    LAYER Metal4 ;
    RECT 452.68 151.795 453.84 160.395 ;
    LAYER Metal4 ;
    RECT 458.08 151.795 459.24 160.395 ;
    LAYER Metal4 ;
    RECT 460.04 151.795 461.2 160.395 ;
    LAYER Metal4 ;
    RECT 465.44 151.795 466.6 160.395 ;
    LAYER Metal4 ;
    RECT 467.4 151.795 468.56 160.395 ;
    LAYER Metal4 ;
    RECT 472.8 151.795 473.96 160.395 ;
    LAYER Metal4 ;
    RECT 474.76 151.795 475.92 160.395 ;
    LAYER Metal4 ;
    RECT 480.16 151.795 481.32 160.395 ;
    LAYER Metal4 ;
    RECT 482.12 151.795 483.28 160.395 ;
    LAYER Metal4 ;
    RECT 487.52 151.795 488.68 160.395 ;
    LAYER Metal4 ;
    RECT 489.48 151.795 490.64 160.395 ;
    LAYER Metal4 ;
    RECT 494.88 151.795 496.04 160.395 ;
    LAYER Metal4 ;
    RECT 496.84 151.795 498 160.395 ;
    LAYER Metal4 ;
    RECT 502.24 151.795 503.4 160.395 ;
    LAYER Metal4 ;
    RECT 504.2 151.795 505.36 160.395 ;
    LAYER Metal4 ;
    RECT 509.6 151.795 510.76 160.395 ;
    LAYER Metal4 ;
    RECT 511.51 151.795 512.61 160.395 ;
    LAYER Metal4 ;
    RECT 513.36 151.795 514.52 160.395 ;
    LAYER Metal4 ;
    RECT 518.76 151.795 519.92 160.395 ;
    LAYER Metal4 ;
    RECT 520.72 151.795 521.88 160.395 ;
    LAYER Metal4 ;
    RECT 526.12 151.795 527.28 160.395 ;
    LAYER Metal4 ;
    RECT 528.08 151.795 529.24 160.395 ;
    LAYER Metal4 ;
    RECT 533.48 151.795 534.64 160.395 ;
    LAYER Metal4 ;
    RECT 535.44 151.795 536.6 160.395 ;
    LAYER Metal4 ;
    RECT 540.84 151.795 542 160.395 ;
    LAYER Metal4 ;
    RECT 542.8 151.795 543.96 160.395 ;
    LAYER Metal4 ;
    RECT 548.2 151.795 549.36 160.395 ;
    LAYER Metal4 ;
    RECT 550.16 151.795 551.32 160.395 ;
    LAYER Metal4 ;
    RECT 555.56 151.795 556.72 160.395 ;
    LAYER Metal4 ;
    RECT 557.52 151.795 558.68 160.395 ;
    LAYER Metal4 ;
    RECT 562.92 151.795 564.08 160.395 ;
    LAYER Metal4 ;
    RECT 564.88 151.795 566.04 160.395 ;
    LAYER Metal4 ;
    RECT 570.28 151.795 571.44 160.395 ;
    LAYER Metal4 ;
    RECT 572.12 151.795 573.4 160.395 ;
    LAYER Metal4 ;
    RECT 19.58 17.2 20.78 8.6 ;
    LAYER Metal4 ;
    RECT 21.48 17.2 22.48 8.6 ;
    LAYER Metal4 ;
    RECT 27.78 17.2 30.9 8.6 ;
    LAYER Metal4 ;
    RECT 36.2 17.2 37.2 8.6 ;
    LAYER Metal4 ;
    RECT 43.1 17.2 44.32 8.6 ;
    LAYER Metal4 ;
    RECT 50.82 17.2 52.02 8.6 ;
    LAYER Metal4 ;
    RECT 58.52 17.2 59.74 8.6 ;
    LAYER Metal4 ;
    RECT 65.64 17.2 66.64 8.6 ;
    LAYER Metal4 ;
    RECT 71.94 17.2 75.06 8.6 ;
    LAYER Metal4 ;
    RECT 80.36 17.2 81.36 8.6 ;
    LAYER Metal4 ;
    RECT 82.16 17.2 83.16 8.6 ;
    LAYER Metal4 ;
    RECT 88.46 17.2 91.58 8.6 ;
    LAYER Metal4 ;
    RECT 96.88 17.2 97.88 8.6 ;
    LAYER Metal4 ;
    RECT 103.78 17.2 105 8.6 ;
    LAYER Metal4 ;
    RECT 111.5 17.2 112.7 8.6 ;
    LAYER Metal4 ;
    RECT 119.2 17.2 120.42 8.6 ;
    LAYER Metal4 ;
    RECT 126.32 17.2 127.32 8.6 ;
    LAYER Metal4 ;
    RECT 132.62 17.2 135.74 8.6 ;
    LAYER Metal4 ;
    RECT 141.04 17.2 142.04 8.6 ;
    LAYER Metal4 ;
    RECT 142.84 17.2 143.84 8.6 ;
    LAYER Metal4 ;
    RECT 149.14 17.2 152.26 8.6 ;
    LAYER Metal4 ;
    RECT 157.56 17.2 158.56 8.6 ;
    LAYER Metal4 ;
    RECT 164.46 17.2 165.68 8.6 ;
    LAYER Metal4 ;
    RECT 172.18 17.2 173.38 8.6 ;
    LAYER Metal4 ;
    RECT 179.88 17.2 181.1 8.6 ;
    LAYER Metal4 ;
    RECT 187 17.2 188 8.6 ;
    LAYER Metal4 ;
    RECT 193.3 17.2 196.42 8.6 ;
    LAYER Metal4 ;
    RECT 201.72 17.2 202.72 8.6 ;
    LAYER Metal4 ;
    RECT 203.52 17.2 204.52 8.6 ;
    LAYER Metal4 ;
    RECT 209.82 17.2 212.94 8.6 ;
    LAYER Metal4 ;
    RECT 218.24 17.2 219.24 8.6 ;
    LAYER Metal4 ;
    RECT 225.14 17.2 226.36 8.6 ;
    LAYER Metal4 ;
    RECT 232.86 17.2 234.06 8.6 ;
    LAYER Metal4 ;
    RECT 240.56 17.2 241.78 8.6 ;
    LAYER Metal4 ;
    RECT 247.68 17.2 248.68 8.6 ;
    LAYER Metal4 ;
    RECT 253.98 17.2 257.1 8.6 ;
    LAYER Metal4 ;
    RECT 262.4 17.2 263.4 8.6 ;
    LAYER Metal4 ;
    RECT 264.2 17.2 265.2 8.6 ;
    LAYER Metal4 ;
    RECT 265.91 17.2 267.51 8.6 ;
    LAYER Metal4 ;
    RECT 268.28 17.2 269.92 8.6 ;
    LAYER Metal4 ;
    RECT 277.08 17.2 278.72 8.6 ;
    LAYER Metal4 ;
    RECT 285.88 17.2 287.52 8.6 ;
    LAYER Metal4 ;
    RECT 294.68 17.2 296.32 8.6 ;
    LAYER Metal4 ;
    RECT 303.48 17.2 305.12 8.6 ;
    LAYER Metal4 ;
    RECT 312.96 17.2 313.82 8.6 ;
    LAYER Metal4 ;
    RECT 318.72 17.2 319.58 8.6 ;
    LAYER Metal4 ;
    RECT 324.48 17.2 325.34 8.6 ;
    LAYER Metal4 ;
    RECT 327.37 17.2 328.35 8.6 ;
    LAYER Metal4 ;
    RECT 330.42 17.2 331.42 8.6 ;
    LAYER Metal4 ;
    RECT 336.72 17.2 339.84 8.6 ;
    LAYER Metal4 ;
    RECT 345.14 17.2 346.14 8.6 ;
    LAYER Metal4 ;
    RECT 352.04 17.2 353.26 8.6 ;
    LAYER Metal4 ;
    RECT 359.76 17.2 360.96 8.6 ;
    LAYER Metal4 ;
    RECT 367.46 17.2 368.68 8.6 ;
    LAYER Metal4 ;
    RECT 374.58 17.2 375.58 8.6 ;
    LAYER Metal4 ;
    RECT 380.88 17.2 384 8.6 ;
    LAYER Metal4 ;
    RECT 389.3 17.2 390.3 8.6 ;
    LAYER Metal4 ;
    RECT 391.1 17.2 392.1 8.6 ;
    LAYER Metal4 ;
    RECT 397.4 17.2 400.52 8.6 ;
    LAYER Metal4 ;
    RECT 405.82 17.2 406.82 8.6 ;
    LAYER Metal4 ;
    RECT 412.72 17.2 413.94 8.6 ;
    LAYER Metal4 ;
    RECT 420.44 17.2 421.64 8.6 ;
    LAYER Metal4 ;
    RECT 428.14 17.2 429.36 8.6 ;
    LAYER Metal4 ;
    RECT 435.26 17.2 436.26 8.6 ;
    LAYER Metal4 ;
    RECT 441.56 17.2 444.68 8.6 ;
    LAYER Metal4 ;
    RECT 449.98 17.2 450.98 8.6 ;
    LAYER Metal4 ;
    RECT 451.78 17.2 452.78 8.6 ;
    LAYER Metal4 ;
    RECT 458.08 17.2 461.2 8.6 ;
    LAYER Metal4 ;
    RECT 466.5 17.2 467.5 8.6 ;
    LAYER Metal4 ;
    RECT 473.4 17.2 474.62 8.6 ;
    LAYER Metal4 ;
    RECT 481.12 17.2 482.32 8.6 ;
    LAYER Metal4 ;
    RECT 488.82 17.2 490.04 8.6 ;
    LAYER Metal4 ;
    RECT 495.94 17.2 496.94 8.6 ;
    LAYER Metal4 ;
    RECT 502.24 17.2 505.36 8.6 ;
    LAYER Metal4 ;
    RECT 510.66 17.2 511.66 8.6 ;
    LAYER Metal4 ;
    RECT 512.46 17.2 513.46 8.6 ;
    LAYER Metal4 ;
    RECT 518.76 17.2 521.88 8.6 ;
    LAYER Metal4 ;
    RECT 527.18 17.2 528.18 8.6 ;
    LAYER Metal4 ;
    RECT 534.08 17.2 535.3 8.6 ;
    LAYER Metal4 ;
    RECT 541.8 17.2 543 8.6 ;
    LAYER Metal4 ;
    RECT 549.5 17.2 550.72 8.6 ;
    LAYER Metal4 ;
    RECT 556.62 17.2 557.62 8.6 ;
    LAYER Metal4 ;
    RECT 562.92 17.2 566.04 8.6 ;
    LAYER Metal4 ;
    RECT 571.34 17.2 572.34 8.6 ;
    LAYER Metal4 ;
    RECT 573.04 17.2 574.24 8.6 ;
    LAYER Metal3 ;
    RECT 576.62 28.715 585.22 30.115 ;
    LAYER Metal3 ;
    RECT 576.62 54.775 585.22 57.275 ;
    LAYER Metal3 ;
    RECT 576.62 63.17 585.22 67.97 ;
    LAYER Metal3 ;
    RECT 576.62 74.265 585.22 74.865 ;
    LAYER Metal3 ;
    RECT 576.62 87.105 585.22 89.105 ;
    LAYER Metal3 ;
    RECT 576.62 121.065 585.22 121.965 ;
    LAYER Metal3 ;
    RECT 576.62 126.125 585.22 127.025 ;
    LAYER Metal3 ;
    RECT 576.62 131.185 585.22 132.085 ;
    LAYER Metal3 ;
    RECT 576.62 136.245 585.22 137.145 ;
    LAYER Metal3 ;
    RECT 576.62 141.305 585.22 142.205 ;
    LAYER Metal3 ;
    RECT 576.62 146.365 585.22 147.265 ;
    LAYER Metal3 ;
    RECT 576.62 149.815 585.22 150.715 ;
    LAYER Metal3 ;
    RECT 17.2 28.715 8.6 30.115 ;
    LAYER Metal3 ;
    RECT 17.2 54.775 8.6 57.275 ;
    LAYER Metal3 ;
    RECT 17.2 63.17 8.6 67.97 ;
    LAYER Metal3 ;
    RECT 17.2 74.265 8.6 74.865 ;
    LAYER Metal3 ;
    RECT 17.2 87.105 8.6 89.105 ;
    LAYER Metal3 ;
    RECT 17.2 121.065 8.6 121.965 ;
    LAYER Metal3 ;
    RECT 17.2 126.125 8.6 127.025 ;
    LAYER Metal3 ;
    RECT 17.2 131.185 8.6 132.085 ;
    LAYER Metal3 ;
    RECT 17.2 136.245 8.6 137.145 ;
    LAYER Metal3 ;
    RECT 17.2 141.305 8.6 142.205 ;
    LAYER Metal3 ;
    RECT 17.2 146.365 8.6 147.265 ;
    LAYER Metal3 ;
    RECT 17.2 149.815 8.6 150.715 ;
    LAYER Via34 ;
    RECT 18.77 161.225 19.55 168.765 ;
    LAYER Via34 ;
    RECT 24.29 161.225 25.07 168.765 ;
    LAYER Via34 ;
    RECT 26.25 161.225 27.03 168.765 ;
    LAYER Via34 ;
    RECT 31.65 161.225 32.43 168.765 ;
    LAYER Via34 ;
    RECT 33.61 161.225 34.39 168.765 ;
    LAYER Via34 ;
    RECT 39.01 161.225 39.79 168.765 ;
    LAYER Via34 ;
    RECT 40.97 161.225 41.75 168.765 ;
    LAYER Via34 ;
    RECT 46.37 161.225 47.15 168.765 ;
    LAYER Via34 ;
    RECT 48.33 161.225 49.11 168.765 ;
    LAYER Via34 ;
    RECT 53.73 161.225 54.51 168.765 ;
    LAYER Via34 ;
    RECT 55.69 161.225 56.47 168.765 ;
    LAYER Via34 ;
    RECT 61.09 161.225 61.87 168.765 ;
    LAYER Via34 ;
    RECT 63.05 161.225 63.83 168.765 ;
    LAYER Via34 ;
    RECT 68.45 161.225 69.23 168.765 ;
    LAYER Via34 ;
    RECT 70.41 161.225 71.19 168.765 ;
    LAYER Via34 ;
    RECT 75.81 161.225 76.59 168.765 ;
    LAYER Via34 ;
    RECT 77.77 161.225 78.55 168.765 ;
    LAYER Via34 ;
    RECT 84.97 161.225 85.75 168.765 ;
    LAYER Via34 ;
    RECT 86.93 161.225 87.71 168.765 ;
    LAYER Via34 ;
    RECT 92.33 161.225 93.11 168.765 ;
    LAYER Via34 ;
    RECT 94.29 161.225 95.07 168.765 ;
    LAYER Via34 ;
    RECT 99.69 161.225 100.47 168.765 ;
    LAYER Via34 ;
    RECT 101.65 161.225 102.43 168.765 ;
    LAYER Via34 ;
    RECT 107.05 161.225 107.83 168.765 ;
    LAYER Via34 ;
    RECT 109.01 161.225 109.79 168.765 ;
    LAYER Via34 ;
    RECT 114.41 161.225 115.19 168.765 ;
    LAYER Via34 ;
    RECT 116.37 161.225 117.15 168.765 ;
    LAYER Via34 ;
    RECT 121.77 161.225 122.55 168.765 ;
    LAYER Via34 ;
    RECT 123.73 161.225 124.51 168.765 ;
    LAYER Via34 ;
    RECT 129.13 161.225 129.91 168.765 ;
    LAYER Via34 ;
    RECT 131.09 161.225 131.87 168.765 ;
    LAYER Via34 ;
    RECT 136.49 161.225 137.27 168.765 ;
    LAYER Via34 ;
    RECT 138.45 161.225 139.23 168.765 ;
    LAYER Via34 ;
    RECT 145.65 161.225 146.43 168.765 ;
    LAYER Via34 ;
    RECT 147.61 161.225 148.39 168.765 ;
    LAYER Via34 ;
    RECT 153.01 161.225 153.79 168.765 ;
    LAYER Via34 ;
    RECT 154.97 161.225 155.75 168.765 ;
    LAYER Via34 ;
    RECT 160.37 161.225 161.15 168.765 ;
    LAYER Via34 ;
    RECT 162.33 161.225 163.11 168.765 ;
    LAYER Via34 ;
    RECT 167.73 161.225 168.51 168.765 ;
    LAYER Via34 ;
    RECT 169.69 161.225 170.47 168.765 ;
    LAYER Via34 ;
    RECT 175.09 161.225 175.87 168.765 ;
    LAYER Via34 ;
    RECT 177.05 161.225 177.83 168.765 ;
    LAYER Via34 ;
    RECT 182.45 161.225 183.23 168.765 ;
    LAYER Via34 ;
    RECT 184.41 161.225 185.19 168.765 ;
    LAYER Via34 ;
    RECT 189.81 161.225 190.59 168.765 ;
    LAYER Via34 ;
    RECT 191.77 161.225 192.55 168.765 ;
    LAYER Via34 ;
    RECT 197.17 161.225 197.95 168.765 ;
    LAYER Via34 ;
    RECT 199.13 161.225 199.91 168.765 ;
    LAYER Via34 ;
    RECT 206.33 161.225 207.11 168.765 ;
    LAYER Via34 ;
    RECT 208.29 161.225 209.07 168.765 ;
    LAYER Via34 ;
    RECT 213.69 161.225 214.47 168.765 ;
    LAYER Via34 ;
    RECT 215.65 161.225 216.43 168.765 ;
    LAYER Via34 ;
    RECT 221.05 161.225 221.83 168.765 ;
    LAYER Via34 ;
    RECT 223.01 161.225 223.79 168.765 ;
    LAYER Via34 ;
    RECT 228.41 161.225 229.19 168.765 ;
    LAYER Via34 ;
    RECT 230.37 161.225 231.15 168.765 ;
    LAYER Via34 ;
    RECT 235.77 161.225 236.55 168.765 ;
    LAYER Via34 ;
    RECT 237.73 161.225 238.51 168.765 ;
    LAYER Via34 ;
    RECT 243.13 161.225 243.91 168.765 ;
    LAYER Via34 ;
    RECT 245.09 161.225 245.87 168.765 ;
    LAYER Via34 ;
    RECT 250.49 161.225 251.27 168.765 ;
    LAYER Via34 ;
    RECT 252.45 161.225 253.23 168.765 ;
    LAYER Via34 ;
    RECT 257.85 161.225 258.63 168.765 ;
    LAYER Via34 ;
    RECT 259.81 161.225 260.59 168.765 ;
    LAYER Via34 ;
    RECT 265.15 161.225 266.45 168.765 ;
    LAYER Via34 ;
    RECT 269.55 161.225 270.85 168.765 ;
    LAYER Via34 ;
    RECT 273.95 161.225 275.25 168.765 ;
    LAYER Via34 ;
    RECT 278.35 161.225 279.65 168.765 ;
    LAYER Via34 ;
    RECT 282.75 161.225 284.05 168.765 ;
    LAYER Via34 ;
    RECT 287.15 161.225 288.45 168.765 ;
    LAYER Via34 ;
    RECT 291.55 161.225 292.85 168.765 ;
    LAYER Via34 ;
    RECT 295.95 161.225 297.25 168.765 ;
    LAYER Via34 ;
    RECT 300.35 161.225 301.65 168.765 ;
    LAYER Via34 ;
    RECT 304.75 161.225 306.05 168.765 ;
    LAYER Via34 ;
    RECT 310.53 161.225 311.31 168.765 ;
    LAYER Via34 ;
    RECT 315.36 161.225 317.18 168.765 ;
    LAYER Via34 ;
    RECT 321.12 161.225 322.94 168.765 ;
    LAYER Via34 ;
    RECT 325.97 161.225 326.75 168.765 ;
    LAYER Via34 ;
    RECT 329.37 161.225 330.67 168.765 ;
    LAYER Via34 ;
    RECT 333.23 161.225 334.01 168.765 ;
    LAYER Via34 ;
    RECT 335.19 161.225 335.97 168.765 ;
    LAYER Via34 ;
    RECT 340.59 161.225 341.37 168.765 ;
    LAYER Via34 ;
    RECT 342.55 161.225 343.33 168.765 ;
    LAYER Via34 ;
    RECT 347.95 161.225 348.73 168.765 ;
    LAYER Via34 ;
    RECT 349.91 161.225 350.69 168.765 ;
    LAYER Via34 ;
    RECT 355.31 161.225 356.09 168.765 ;
    LAYER Via34 ;
    RECT 357.27 161.225 358.05 168.765 ;
    LAYER Via34 ;
    RECT 362.67 161.225 363.45 168.765 ;
    LAYER Via34 ;
    RECT 364.63 161.225 365.41 168.765 ;
    LAYER Via34 ;
    RECT 370.03 161.225 370.81 168.765 ;
    LAYER Via34 ;
    RECT 371.99 161.225 372.77 168.765 ;
    LAYER Via34 ;
    RECT 377.39 161.225 378.17 168.765 ;
    LAYER Via34 ;
    RECT 379.35 161.225 380.13 168.765 ;
    LAYER Via34 ;
    RECT 384.75 161.225 385.53 168.765 ;
    LAYER Via34 ;
    RECT 386.71 161.225 387.49 168.765 ;
    LAYER Via34 ;
    RECT 393.91 161.225 394.69 168.765 ;
    LAYER Via34 ;
    RECT 395.87 161.225 396.65 168.765 ;
    LAYER Via34 ;
    RECT 401.27 161.225 402.05 168.765 ;
    LAYER Via34 ;
    RECT 403.23 161.225 404.01 168.765 ;
    LAYER Via34 ;
    RECT 408.63 161.225 409.41 168.765 ;
    LAYER Via34 ;
    RECT 410.59 161.225 411.37 168.765 ;
    LAYER Via34 ;
    RECT 415.99 161.225 416.77 168.765 ;
    LAYER Via34 ;
    RECT 417.95 161.225 418.73 168.765 ;
    LAYER Via34 ;
    RECT 423.35 161.225 424.13 168.765 ;
    LAYER Via34 ;
    RECT 425.31 161.225 426.09 168.765 ;
    LAYER Via34 ;
    RECT 430.71 161.225 431.49 168.765 ;
    LAYER Via34 ;
    RECT 432.67 161.225 433.45 168.765 ;
    LAYER Via34 ;
    RECT 438.07 161.225 438.85 168.765 ;
    LAYER Via34 ;
    RECT 440.03 161.225 440.81 168.765 ;
    LAYER Via34 ;
    RECT 445.43 161.225 446.21 168.765 ;
    LAYER Via34 ;
    RECT 447.39 161.225 448.17 168.765 ;
    LAYER Via34 ;
    RECT 454.59 161.225 455.37 168.765 ;
    LAYER Via34 ;
    RECT 456.55 161.225 457.33 168.765 ;
    LAYER Via34 ;
    RECT 461.95 161.225 462.73 168.765 ;
    LAYER Via34 ;
    RECT 463.91 161.225 464.69 168.765 ;
    LAYER Via34 ;
    RECT 469.31 161.225 470.09 168.765 ;
    LAYER Via34 ;
    RECT 471.27 161.225 472.05 168.765 ;
    LAYER Via34 ;
    RECT 476.67 161.225 477.45 168.765 ;
    LAYER Via34 ;
    RECT 478.63 161.225 479.41 168.765 ;
    LAYER Via34 ;
    RECT 484.03 161.225 484.81 168.765 ;
    LAYER Via34 ;
    RECT 485.99 161.225 486.77 168.765 ;
    LAYER Via34 ;
    RECT 491.39 161.225 492.17 168.765 ;
    LAYER Via34 ;
    RECT 493.35 161.225 494.13 168.765 ;
    LAYER Via34 ;
    RECT 498.75 161.225 499.53 168.765 ;
    LAYER Via34 ;
    RECT 500.71 161.225 501.49 168.765 ;
    LAYER Via34 ;
    RECT 506.11 161.225 506.89 168.765 ;
    LAYER Via34 ;
    RECT 508.07 161.225 508.85 168.765 ;
    LAYER Via34 ;
    RECT 515.27 161.225 516.05 168.765 ;
    LAYER Via34 ;
    RECT 517.23 161.225 518.01 168.765 ;
    LAYER Via34 ;
    RECT 522.63 161.225 523.41 168.765 ;
    LAYER Via34 ;
    RECT 524.59 161.225 525.37 168.765 ;
    LAYER Via34 ;
    RECT 529.99 161.225 530.77 168.765 ;
    LAYER Via34 ;
    RECT 531.95 161.225 532.73 168.765 ;
    LAYER Via34 ;
    RECT 537.35 161.225 538.13 168.765 ;
    LAYER Via34 ;
    RECT 539.31 161.225 540.09 168.765 ;
    LAYER Via34 ;
    RECT 544.71 161.225 545.49 168.765 ;
    LAYER Via34 ;
    RECT 546.67 161.225 547.45 168.765 ;
    LAYER Via34 ;
    RECT 552.07 161.225 552.85 168.765 ;
    LAYER Via34 ;
    RECT 554.03 161.225 554.81 168.765 ;
    LAYER Via34 ;
    RECT 559.43 161.225 560.21 168.765 ;
    LAYER Via34 ;
    RECT 561.39 161.225 562.17 168.765 ;
    LAYER Via34 ;
    RECT 566.79 161.225 567.57 168.765 ;
    LAYER Via34 ;
    RECT 568.75 161.225 569.53 168.765 ;
    LAYER Via34 ;
    RECT 574.27 161.225 575.05 168.765 ;
    LAYER Via34 ;
    RECT 18.18 0.23 18.96 7.77 ;
    LAYER Via34 ;
    RECT 24.23 0.23 27.09 7.77 ;
    LAYER Via34 ;
    RECT 31.59 0.23 34.45 7.77 ;
    LAYER Via34 ;
    RECT 38.46 0.23 39.24 7.77 ;
    LAYER Via34 ;
    RECT 47.3 0.23 49.12 7.77 ;
    LAYER Via34 ;
    RECT 53.72 0.23 55.54 7.77 ;
    LAYER Via34 ;
    RECT 63.6 0.23 64.38 7.77 ;
    LAYER Via34 ;
    RECT 68.39 0.23 71.25 7.77 ;
    LAYER Via34 ;
    RECT 75.75 0.23 78.61 7.77 ;
    LAYER Via34 ;
    RECT 84.91 0.23 87.77 7.77 ;
    LAYER Via34 ;
    RECT 92.27 0.23 95.13 7.77 ;
    LAYER Via34 ;
    RECT 99.14 0.23 99.92 7.77 ;
    LAYER Via34 ;
    RECT 107.98 0.23 109.8 7.77 ;
    LAYER Via34 ;
    RECT 114.4 0.23 116.22 7.77 ;
    LAYER Via34 ;
    RECT 124.28 0.23 125.06 7.77 ;
    LAYER Via34 ;
    RECT 129.07 0.23 131.93 7.77 ;
    LAYER Via34 ;
    RECT 136.43 0.23 139.29 7.77 ;
    LAYER Via34 ;
    RECT 145.59 0.23 148.45 7.77 ;
    LAYER Via34 ;
    RECT 152.95 0.23 155.81 7.77 ;
    LAYER Via34 ;
    RECT 159.82 0.23 160.6 7.77 ;
    LAYER Via34 ;
    RECT 168.66 0.23 170.48 7.77 ;
    LAYER Via34 ;
    RECT 175.08 0.23 176.9 7.77 ;
    LAYER Via34 ;
    RECT 184.96 0.23 185.74 7.77 ;
    LAYER Via34 ;
    RECT 189.75 0.23 192.61 7.77 ;
    LAYER Via34 ;
    RECT 197.11 0.23 199.97 7.77 ;
    LAYER Via34 ;
    RECT 206.27 0.23 209.13 7.77 ;
    LAYER Via34 ;
    RECT 213.63 0.23 216.49 7.77 ;
    LAYER Via34 ;
    RECT 220.5 0.23 221.28 7.77 ;
    LAYER Via34 ;
    RECT 229.34 0.23 231.16 7.77 ;
    LAYER Via34 ;
    RECT 235.76 0.23 237.58 7.77 ;
    LAYER Via34 ;
    RECT 245.64 0.23 246.42 7.77 ;
    LAYER Via34 ;
    RECT 250.43 0.23 253.29 7.77 ;
    LAYER Via34 ;
    RECT 257.79 0.23 260.65 7.77 ;
    LAYER Via34 ;
    RECT 270.79 0.23 274.17 7.77 ;
    LAYER Via34 ;
    RECT 281.65 0.23 282.95 7.77 ;
    LAYER Via34 ;
    RECT 288.39 0.23 291.77 7.77 ;
    LAYER Via34 ;
    RECT 299.25 0.23 300.55 7.77 ;
    LAYER Via34 ;
    RECT 308.57 0.23 308.83 7.77 ;
    LAYER Via34 ;
    RECT 310.12 0.23 310.9 7.77 ;
    LAYER Via34 ;
    RECT 316.14 0.23 316.4 7.77 ;
    LAYER Via34 ;
    RECT 321.9 0.23 322.16 7.77 ;
    LAYER Via34 ;
    RECT 333.17 0.23 336.03 7.77 ;
    LAYER Via34 ;
    RECT 340.53 0.23 343.39 7.77 ;
    LAYER Via34 ;
    RECT 347.4 0.23 348.18 7.77 ;
    LAYER Via34 ;
    RECT 356.24 0.23 358.06 7.77 ;
    LAYER Via34 ;
    RECT 362.66 0.23 364.48 7.77 ;
    LAYER Via34 ;
    RECT 372.54 0.23 373.32 7.77 ;
    LAYER Via34 ;
    RECT 377.33 0.23 380.19 7.77 ;
    LAYER Via34 ;
    RECT 384.69 0.23 387.55 7.77 ;
    LAYER Via34 ;
    RECT 393.85 0.23 396.71 7.77 ;
    LAYER Via34 ;
    RECT 401.21 0.23 404.07 7.77 ;
    LAYER Via34 ;
    RECT 408.08 0.23 408.86 7.77 ;
    LAYER Via34 ;
    RECT 416.92 0.23 418.74 7.77 ;
    LAYER Via34 ;
    RECT 423.34 0.23 425.16 7.77 ;
    LAYER Via34 ;
    RECT 433.22 0.23 434 7.77 ;
    LAYER Via34 ;
    RECT 438.01 0.23 440.87 7.77 ;
    LAYER Via34 ;
    RECT 445.37 0.23 448.23 7.77 ;
    LAYER Via34 ;
    RECT 454.53 0.23 457.39 7.77 ;
    LAYER Via34 ;
    RECT 461.89 0.23 464.75 7.77 ;
    LAYER Via34 ;
    RECT 468.76 0.23 469.54 7.77 ;
    LAYER Via34 ;
    RECT 477.6 0.23 479.42 7.77 ;
    LAYER Via34 ;
    RECT 484.02 0.23 485.84 7.77 ;
    LAYER Via34 ;
    RECT 493.9 0.23 494.68 7.77 ;
    LAYER Via34 ;
    RECT 498.69 0.23 501.55 7.77 ;
    LAYER Via34 ;
    RECT 506.05 0.23 508.91 7.77 ;
    LAYER Via34 ;
    RECT 515.21 0.23 518.07 7.77 ;
    LAYER Via34 ;
    RECT 522.57 0.23 525.43 7.77 ;
    LAYER Via34 ;
    RECT 529.44 0.23 530.22 7.77 ;
    LAYER Via34 ;
    RECT 538.28 0.23 540.1 7.77 ;
    LAYER Via34 ;
    RECT 544.7 0.23 546.52 7.77 ;
    LAYER Via34 ;
    RECT 554.58 0.23 555.36 7.77 ;
    LAYER Via34 ;
    RECT 559.37 0.23 562.23 7.77 ;
    LAYER Via34 ;
    RECT 566.73 0.23 569.59 7.77 ;
    LAYER Via34 ;
    RECT 574.86 0.23 575.64 7.77 ;
    LAYER Via34 ;
    RECT 586.05 22.33 593.59 23.11 ;
    LAYER Via34 ;
    RECT 586.05 35.2 593.59 35.98 ;
    LAYER Via34 ;
    RECT 586.05 48.415 593.59 48.675 ;
    LAYER Via34 ;
    RECT 586.05 52.665 593.59 53.445 ;
    LAYER Via34 ;
    RECT 586.05 73.375 593.59 73.635 ;
    LAYER Via34 ;
    RECT 586.05 82.835 593.59 84.135 ;
    LAYER Via34 ;
    RECT 586.05 90.41 593.59 94.31 ;
    LAYER Via34 ;
    RECT 586.05 95.38 593.59 103.44 ;
    LAYER Via34 ;
    RECT 586.05 106.035 593.59 109.415 ;
    LAYER Via34 ;
    RECT 586.05 110.5 593.59 113.88 ;
    LAYER Via34 ;
    RECT 586.05 123.655 593.59 124.435 ;
    LAYER Via34 ;
    RECT 586.05 128.715 593.59 129.495 ;
    LAYER Via34 ;
    RECT 586.05 133.775 593.59 134.555 ;
    LAYER Via34 ;
    RECT 586.05 138.835 593.59 139.615 ;
    LAYER Via34 ;
    RECT 586.05 144.165 593.59 144.945 ;
    LAYER Via34 ;
    RECT 586.05 148.065 593.59 148.845 ;
    LAYER Via34 ;
    RECT 0.23 22.33 7.77 23.11 ;
    LAYER Via34 ;
    RECT 0.23 35.2 7.77 35.98 ;
    LAYER Via34 ;
    RECT 0.23 48.415 7.77 48.675 ;
    LAYER Via34 ;
    RECT 0.23 52.665 7.77 53.445 ;
    LAYER Via34 ;
    RECT 0.23 73.375 7.77 73.635 ;
    LAYER Via34 ;
    RECT 0.23 82.835 7.77 84.135 ;
    LAYER Via34 ;
    RECT 0.23 90.41 7.77 94.31 ;
    LAYER Via34 ;
    RECT 0.23 95.38 7.77 103.44 ;
    LAYER Via34 ;
    RECT 0.23 106.035 7.77 109.415 ;
    LAYER Via34 ;
    RECT 0.23 110.5 7.77 113.88 ;
    LAYER Via34 ;
    RECT 0.23 123.655 7.77 124.435 ;
    LAYER Via34 ;
    RECT 0.23 128.715 7.77 129.495 ;
    LAYER Via34 ;
    RECT 0.23 133.775 7.77 134.555 ;
    LAYER Via34 ;
    RECT 0.23 138.835 7.77 139.615 ;
    LAYER Via34 ;
    RECT 0.23 144.165 7.77 144.945 ;
    LAYER Via34 ;
    RECT 0.23 148.065 7.77 148.845 ;
    LAYER Via34 ;
    RECT 20.67 152.625 21.45 160.165 ;
    LAYER Via34 ;
    RECT 22.57 152.625 23.35 160.165 ;
    LAYER Via34 ;
    RECT 27.97 152.625 28.75 160.165 ;
    LAYER Via34 ;
    RECT 29.93 152.625 30.71 160.165 ;
    LAYER Via34 ;
    RECT 35.33 152.625 36.11 160.165 ;
    LAYER Via34 ;
    RECT 37.29 152.625 38.07 160.165 ;
    LAYER Via34 ;
    RECT 42.69 152.625 43.47 160.165 ;
    LAYER Via34 ;
    RECT 44.65 152.625 45.43 160.165 ;
    LAYER Via34 ;
    RECT 50.05 152.625 50.83 160.165 ;
    LAYER Via34 ;
    RECT 52.01 152.625 52.79 160.165 ;
    LAYER Via34 ;
    RECT 57.41 152.625 58.19 160.165 ;
    LAYER Via34 ;
    RECT 59.37 152.625 60.15 160.165 ;
    LAYER Via34 ;
    RECT 64.77 152.625 65.55 160.165 ;
    LAYER Via34 ;
    RECT 66.73 152.625 67.51 160.165 ;
    LAYER Via34 ;
    RECT 72.13 152.625 72.91 160.165 ;
    LAYER Via34 ;
    RECT 74.09 152.625 74.87 160.165 ;
    LAYER Via34 ;
    RECT 79.49 152.625 80.27 160.165 ;
    LAYER Via34 ;
    RECT 81.37 152.625 82.15 160.165 ;
    LAYER Via34 ;
    RECT 83.25 152.625 84.03 160.165 ;
    LAYER Via34 ;
    RECT 88.65 152.625 89.43 160.165 ;
    LAYER Via34 ;
    RECT 90.61 152.625 91.39 160.165 ;
    LAYER Via34 ;
    RECT 96.01 152.625 96.79 160.165 ;
    LAYER Via34 ;
    RECT 97.97 152.625 98.75 160.165 ;
    LAYER Via34 ;
    RECT 103.37 152.625 104.15 160.165 ;
    LAYER Via34 ;
    RECT 105.33 152.625 106.11 160.165 ;
    LAYER Via34 ;
    RECT 110.73 152.625 111.51 160.165 ;
    LAYER Via34 ;
    RECT 112.69 152.625 113.47 160.165 ;
    LAYER Via34 ;
    RECT 118.09 152.625 118.87 160.165 ;
    LAYER Via34 ;
    RECT 120.05 152.625 120.83 160.165 ;
    LAYER Via34 ;
    RECT 125.45 152.625 126.23 160.165 ;
    LAYER Via34 ;
    RECT 127.41 152.625 128.19 160.165 ;
    LAYER Via34 ;
    RECT 132.81 152.625 133.59 160.165 ;
    LAYER Via34 ;
    RECT 134.77 152.625 135.55 160.165 ;
    LAYER Via34 ;
    RECT 140.17 152.625 140.95 160.165 ;
    LAYER Via34 ;
    RECT 142.05 152.625 142.83 160.165 ;
    LAYER Via34 ;
    RECT 143.93 152.625 144.71 160.165 ;
    LAYER Via34 ;
    RECT 149.33 152.625 150.11 160.165 ;
    LAYER Via34 ;
    RECT 151.29 152.625 152.07 160.165 ;
    LAYER Via34 ;
    RECT 156.69 152.625 157.47 160.165 ;
    LAYER Via34 ;
    RECT 158.65 152.625 159.43 160.165 ;
    LAYER Via34 ;
    RECT 164.05 152.625 164.83 160.165 ;
    LAYER Via34 ;
    RECT 166.01 152.625 166.79 160.165 ;
    LAYER Via34 ;
    RECT 171.41 152.625 172.19 160.165 ;
    LAYER Via34 ;
    RECT 173.37 152.625 174.15 160.165 ;
    LAYER Via34 ;
    RECT 178.77 152.625 179.55 160.165 ;
    LAYER Via34 ;
    RECT 180.73 152.625 181.51 160.165 ;
    LAYER Via34 ;
    RECT 186.13 152.625 186.91 160.165 ;
    LAYER Via34 ;
    RECT 188.09 152.625 188.87 160.165 ;
    LAYER Via34 ;
    RECT 193.49 152.625 194.27 160.165 ;
    LAYER Via34 ;
    RECT 195.45 152.625 196.23 160.165 ;
    LAYER Via34 ;
    RECT 200.85 152.625 201.63 160.165 ;
    LAYER Via34 ;
    RECT 202.73 152.625 203.51 160.165 ;
    LAYER Via34 ;
    RECT 204.61 152.625 205.39 160.165 ;
    LAYER Via34 ;
    RECT 210.01 152.625 210.79 160.165 ;
    LAYER Via34 ;
    RECT 211.97 152.625 212.75 160.165 ;
    LAYER Via34 ;
    RECT 217.37 152.625 218.15 160.165 ;
    LAYER Via34 ;
    RECT 219.33 152.625 220.11 160.165 ;
    LAYER Via34 ;
    RECT 224.73 152.625 225.51 160.165 ;
    LAYER Via34 ;
    RECT 226.69 152.625 227.47 160.165 ;
    LAYER Via34 ;
    RECT 232.09 152.625 232.87 160.165 ;
    LAYER Via34 ;
    RECT 234.05 152.625 234.83 160.165 ;
    LAYER Via34 ;
    RECT 239.45 152.625 240.23 160.165 ;
    LAYER Via34 ;
    RECT 241.41 152.625 242.19 160.165 ;
    LAYER Via34 ;
    RECT 246.81 152.625 247.59 160.165 ;
    LAYER Via34 ;
    RECT 248.77 152.625 249.55 160.165 ;
    LAYER Via34 ;
    RECT 254.17 152.625 254.95 160.165 ;
    LAYER Via34 ;
    RECT 256.13 152.625 256.91 160.165 ;
    LAYER Via34 ;
    RECT 261.53 152.625 262.31 160.165 ;
    LAYER Via34 ;
    RECT 263.41 152.625 264.19 160.165 ;
    LAYER Via34 ;
    RECT 267.35 152.625 268.65 160.165 ;
    LAYER Via34 ;
    RECT 271.75 152.625 273.05 160.165 ;
    LAYER Via34 ;
    RECT 276.15 152.625 277.45 160.165 ;
    LAYER Via34 ;
    RECT 280.55 152.625 281.85 160.165 ;
    LAYER Via34 ;
    RECT 284.95 152.625 286.25 160.165 ;
    LAYER Via34 ;
    RECT 289.35 152.625 290.65 160.165 ;
    LAYER Via34 ;
    RECT 293.75 152.625 295.05 160.165 ;
    LAYER Via34 ;
    RECT 298.15 152.625 299.45 160.165 ;
    LAYER Via34 ;
    RECT 302.55 152.625 303.85 160.165 ;
    LAYER Via34 ;
    RECT 306.77 152.625 309.63 160.165 ;
    LAYER Via34 ;
    RECT 312.48 152.625 314.3 160.165 ;
    LAYER Via34 ;
    RECT 318.24 152.625 320.06 160.165 ;
    LAYER Via34 ;
    RECT 324.11 152.625 324.89 160.165 ;
    LAYER Via34 ;
    RECT 327.81 152.625 328.59 160.165 ;
    LAYER Via34 ;
    RECT 331.51 152.625 332.29 160.165 ;
    LAYER Via34 ;
    RECT 336.91 152.625 337.69 160.165 ;
    LAYER Via34 ;
    RECT 338.87 152.625 339.65 160.165 ;
    LAYER Via34 ;
    RECT 344.27 152.625 345.05 160.165 ;
    LAYER Via34 ;
    RECT 346.23 152.625 347.01 160.165 ;
    LAYER Via34 ;
    RECT 351.63 152.625 352.41 160.165 ;
    LAYER Via34 ;
    RECT 353.59 152.625 354.37 160.165 ;
    LAYER Via34 ;
    RECT 358.99 152.625 359.77 160.165 ;
    LAYER Via34 ;
    RECT 360.95 152.625 361.73 160.165 ;
    LAYER Via34 ;
    RECT 366.35 152.625 367.13 160.165 ;
    LAYER Via34 ;
    RECT 368.31 152.625 369.09 160.165 ;
    LAYER Via34 ;
    RECT 373.71 152.625 374.49 160.165 ;
    LAYER Via34 ;
    RECT 375.67 152.625 376.45 160.165 ;
    LAYER Via34 ;
    RECT 381.07 152.625 381.85 160.165 ;
    LAYER Via34 ;
    RECT 383.03 152.625 383.81 160.165 ;
    LAYER Via34 ;
    RECT 388.43 152.625 389.21 160.165 ;
    LAYER Via34 ;
    RECT 390.31 152.625 391.09 160.165 ;
    LAYER Via34 ;
    RECT 392.19 152.625 392.97 160.165 ;
    LAYER Via34 ;
    RECT 397.59 152.625 398.37 160.165 ;
    LAYER Via34 ;
    RECT 399.55 152.625 400.33 160.165 ;
    LAYER Via34 ;
    RECT 404.95 152.625 405.73 160.165 ;
    LAYER Via34 ;
    RECT 406.91 152.625 407.69 160.165 ;
    LAYER Via34 ;
    RECT 412.31 152.625 413.09 160.165 ;
    LAYER Via34 ;
    RECT 414.27 152.625 415.05 160.165 ;
    LAYER Via34 ;
    RECT 419.67 152.625 420.45 160.165 ;
    LAYER Via34 ;
    RECT 421.63 152.625 422.41 160.165 ;
    LAYER Via34 ;
    RECT 427.03 152.625 427.81 160.165 ;
    LAYER Via34 ;
    RECT 428.99 152.625 429.77 160.165 ;
    LAYER Via34 ;
    RECT 434.39 152.625 435.17 160.165 ;
    LAYER Via34 ;
    RECT 436.35 152.625 437.13 160.165 ;
    LAYER Via34 ;
    RECT 441.75 152.625 442.53 160.165 ;
    LAYER Via34 ;
    RECT 443.71 152.625 444.49 160.165 ;
    LAYER Via34 ;
    RECT 449.11 152.625 449.89 160.165 ;
    LAYER Via34 ;
    RECT 450.99 152.625 451.77 160.165 ;
    LAYER Via34 ;
    RECT 452.87 152.625 453.65 160.165 ;
    LAYER Via34 ;
    RECT 458.27 152.625 459.05 160.165 ;
    LAYER Via34 ;
    RECT 460.23 152.625 461.01 160.165 ;
    LAYER Via34 ;
    RECT 465.63 152.625 466.41 160.165 ;
    LAYER Via34 ;
    RECT 467.59 152.625 468.37 160.165 ;
    LAYER Via34 ;
    RECT 472.99 152.625 473.77 160.165 ;
    LAYER Via34 ;
    RECT 474.95 152.625 475.73 160.165 ;
    LAYER Via34 ;
    RECT 480.35 152.625 481.13 160.165 ;
    LAYER Via34 ;
    RECT 482.31 152.625 483.09 160.165 ;
    LAYER Via34 ;
    RECT 487.71 152.625 488.49 160.165 ;
    LAYER Via34 ;
    RECT 489.67 152.625 490.45 160.165 ;
    LAYER Via34 ;
    RECT 495.07 152.625 495.85 160.165 ;
    LAYER Via34 ;
    RECT 497.03 152.625 497.81 160.165 ;
    LAYER Via34 ;
    RECT 502.43 152.625 503.21 160.165 ;
    LAYER Via34 ;
    RECT 504.39 152.625 505.17 160.165 ;
    LAYER Via34 ;
    RECT 509.79 152.625 510.57 160.165 ;
    LAYER Via34 ;
    RECT 511.67 152.625 512.45 160.165 ;
    LAYER Via34 ;
    RECT 513.55 152.625 514.33 160.165 ;
    LAYER Via34 ;
    RECT 518.95 152.625 519.73 160.165 ;
    LAYER Via34 ;
    RECT 520.91 152.625 521.69 160.165 ;
    LAYER Via34 ;
    RECT 526.31 152.625 527.09 160.165 ;
    LAYER Via34 ;
    RECT 528.27 152.625 529.05 160.165 ;
    LAYER Via34 ;
    RECT 533.67 152.625 534.45 160.165 ;
    LAYER Via34 ;
    RECT 535.63 152.625 536.41 160.165 ;
    LAYER Via34 ;
    RECT 541.03 152.625 541.81 160.165 ;
    LAYER Via34 ;
    RECT 542.99 152.625 543.77 160.165 ;
    LAYER Via34 ;
    RECT 548.39 152.625 549.17 160.165 ;
    LAYER Via34 ;
    RECT 550.35 152.625 551.13 160.165 ;
    LAYER Via34 ;
    RECT 555.75 152.625 556.53 160.165 ;
    LAYER Via34 ;
    RECT 557.71 152.625 558.49 160.165 ;
    LAYER Via34 ;
    RECT 563.11 152.625 563.89 160.165 ;
    LAYER Via34 ;
    RECT 565.07 152.625 565.85 160.165 ;
    LAYER Via34 ;
    RECT 570.47 152.625 571.25 160.165 ;
    LAYER Via34 ;
    RECT 572.37 152.625 573.15 160.165 ;
    LAYER Via34 ;
    RECT 19.79 8.83 20.57 16.37 ;
    LAYER Via34 ;
    RECT 21.59 8.83 22.37 16.37 ;
    LAYER Via34 ;
    RECT 27.91 8.83 30.77 16.37 ;
    LAYER Via34 ;
    RECT 36.31 8.83 37.09 16.37 ;
    LAYER Via34 ;
    RECT 43.32 8.83 44.1 16.37 ;
    LAYER Via34 ;
    RECT 51.03 8.83 51.81 16.37 ;
    LAYER Via34 ;
    RECT 58.74 8.83 59.52 16.37 ;
    LAYER Via34 ;
    RECT 65.75 8.83 66.53 16.37 ;
    LAYER Via34 ;
    RECT 72.07 8.83 74.93 16.37 ;
    LAYER Via34 ;
    RECT 80.47 8.83 81.25 16.37 ;
    LAYER Via34 ;
    RECT 82.27 8.83 83.05 16.37 ;
    LAYER Via34 ;
    RECT 88.59 8.83 91.45 16.37 ;
    LAYER Via34 ;
    RECT 96.99 8.83 97.77 16.37 ;
    LAYER Via34 ;
    RECT 104 8.83 104.78 16.37 ;
    LAYER Via34 ;
    RECT 111.71 8.83 112.49 16.37 ;
    LAYER Via34 ;
    RECT 119.42 8.83 120.2 16.37 ;
    LAYER Via34 ;
    RECT 126.43 8.83 127.21 16.37 ;
    LAYER Via34 ;
    RECT 132.75 8.83 135.61 16.37 ;
    LAYER Via34 ;
    RECT 141.15 8.83 141.93 16.37 ;
    LAYER Via34 ;
    RECT 142.95 8.83 143.73 16.37 ;
    LAYER Via34 ;
    RECT 149.27 8.83 152.13 16.37 ;
    LAYER Via34 ;
    RECT 157.67 8.83 158.45 16.37 ;
    LAYER Via34 ;
    RECT 164.68 8.83 165.46 16.37 ;
    LAYER Via34 ;
    RECT 172.39 8.83 173.17 16.37 ;
    LAYER Via34 ;
    RECT 180.1 8.83 180.88 16.37 ;
    LAYER Via34 ;
    RECT 187.11 8.83 187.89 16.37 ;
    LAYER Via34 ;
    RECT 193.43 8.83 196.29 16.37 ;
    LAYER Via34 ;
    RECT 201.83 8.83 202.61 16.37 ;
    LAYER Via34 ;
    RECT 203.63 8.83 204.41 16.37 ;
    LAYER Via34 ;
    RECT 209.95 8.83 212.81 16.37 ;
    LAYER Via34 ;
    RECT 218.35 8.83 219.13 16.37 ;
    LAYER Via34 ;
    RECT 225.36 8.83 226.14 16.37 ;
    LAYER Via34 ;
    RECT 233.07 8.83 233.85 16.37 ;
    LAYER Via34 ;
    RECT 240.78 8.83 241.56 16.37 ;
    LAYER Via34 ;
    RECT 247.79 8.83 248.57 16.37 ;
    LAYER Via34 ;
    RECT 254.11 8.83 256.97 16.37 ;
    LAYER Via34 ;
    RECT 262.51 8.83 263.29 16.37 ;
    LAYER Via34 ;
    RECT 264.31 8.83 265.09 16.37 ;
    LAYER Via34 ;
    RECT 266.06 8.83 267.36 16.37 ;
    LAYER Via34 ;
    RECT 268.45 8.83 269.75 16.37 ;
    LAYER Via34 ;
    RECT 277.25 8.83 278.55 16.37 ;
    LAYER Via34 ;
    RECT 286.05 8.83 287.35 16.37 ;
    LAYER Via34 ;
    RECT 294.85 8.83 296.15 16.37 ;
    LAYER Via34 ;
    RECT 303.65 8.83 304.95 16.37 ;
    LAYER Via34 ;
    RECT 313.26 8.83 313.52 16.37 ;
    LAYER Via34 ;
    RECT 319.02 8.83 319.28 16.37 ;
    LAYER Via34 ;
    RECT 324.78 8.83 325.04 16.37 ;
    LAYER Via34 ;
    RECT 327.47 8.83 328.25 16.37 ;
    LAYER Via34 ;
    RECT 330.53 8.83 331.31 16.37 ;
    LAYER Via34 ;
    RECT 336.85 8.83 339.71 16.37 ;
    LAYER Via34 ;
    RECT 345.25 8.83 346.03 16.37 ;
    LAYER Via34 ;
    RECT 352.26 8.83 353.04 16.37 ;
    LAYER Via34 ;
    RECT 359.97 8.83 360.75 16.37 ;
    LAYER Via34 ;
    RECT 367.68 8.83 368.46 16.37 ;
    LAYER Via34 ;
    RECT 374.69 8.83 375.47 16.37 ;
    LAYER Via34 ;
    RECT 381.01 8.83 383.87 16.37 ;
    LAYER Via34 ;
    RECT 389.41 8.83 390.19 16.37 ;
    LAYER Via34 ;
    RECT 391.21 8.83 391.99 16.37 ;
    LAYER Via34 ;
    RECT 397.53 8.83 400.39 16.37 ;
    LAYER Via34 ;
    RECT 405.93 8.83 406.71 16.37 ;
    LAYER Via34 ;
    RECT 412.94 8.83 413.72 16.37 ;
    LAYER Via34 ;
    RECT 420.65 8.83 421.43 16.37 ;
    LAYER Via34 ;
    RECT 428.36 8.83 429.14 16.37 ;
    LAYER Via34 ;
    RECT 435.37 8.83 436.15 16.37 ;
    LAYER Via34 ;
    RECT 441.69 8.83 444.55 16.37 ;
    LAYER Via34 ;
    RECT 450.09 8.83 450.87 16.37 ;
    LAYER Via34 ;
    RECT 451.89 8.83 452.67 16.37 ;
    LAYER Via34 ;
    RECT 458.21 8.83 461.07 16.37 ;
    LAYER Via34 ;
    RECT 466.61 8.83 467.39 16.37 ;
    LAYER Via34 ;
    RECT 473.62 8.83 474.4 16.37 ;
    LAYER Via34 ;
    RECT 481.33 8.83 482.11 16.37 ;
    LAYER Via34 ;
    RECT 489.04 8.83 489.82 16.37 ;
    LAYER Via34 ;
    RECT 496.05 8.83 496.83 16.37 ;
    LAYER Via34 ;
    RECT 502.37 8.83 505.23 16.37 ;
    LAYER Via34 ;
    RECT 510.77 8.83 511.55 16.37 ;
    LAYER Via34 ;
    RECT 512.57 8.83 513.35 16.37 ;
    LAYER Via34 ;
    RECT 518.89 8.83 521.75 16.37 ;
    LAYER Via34 ;
    RECT 527.29 8.83 528.07 16.37 ;
    LAYER Via34 ;
    RECT 534.3 8.83 535.08 16.37 ;
    LAYER Via34 ;
    RECT 542.01 8.83 542.79 16.37 ;
    LAYER Via34 ;
    RECT 549.72 8.83 550.5 16.37 ;
    LAYER Via34 ;
    RECT 556.73 8.83 557.51 16.37 ;
    LAYER Via34 ;
    RECT 563.05 8.83 565.91 16.37 ;
    LAYER Via34 ;
    RECT 571.45 8.83 572.23 16.37 ;
    LAYER Via34 ;
    RECT 573.25 8.83 574.03 16.37 ;
    LAYER Via34 ;
    RECT 577.45 29.025 584.99 29.805 ;
    LAYER Via34 ;
    RECT 577.45 54.855 584.99 57.195 ;
    LAYER Via34 ;
    RECT 577.45 63.36 584.99 67.78 ;
    LAYER Via34 ;
    RECT 577.45 74.435 584.99 74.695 ;
    LAYER Via34 ;
    RECT 577.45 87.195 584.99 89.015 ;
    LAYER Via34 ;
    RECT 577.45 121.125 584.99 121.905 ;
    LAYER Via34 ;
    RECT 577.45 126.185 584.99 126.965 ;
    LAYER Via34 ;
    RECT 577.45 131.245 584.99 132.025 ;
    LAYER Via34 ;
    RECT 577.45 136.305 584.99 137.085 ;
    LAYER Via34 ;
    RECT 577.45 141.365 584.99 142.145 ;
    LAYER Via34 ;
    RECT 577.45 146.425 584.99 147.205 ;
    LAYER Via34 ;
    RECT 577.45 149.875 584.99 150.655 ;
    LAYER Via34 ;
    RECT 8.83 29.025 16.37 29.805 ;
    LAYER Via34 ;
    RECT 8.83 54.855 16.37 57.195 ;
    LAYER Via34 ;
    RECT 8.83 63.36 16.37 67.78 ;
    LAYER Via34 ;
    RECT 8.83 74.435 16.37 74.695 ;
    LAYER Via34 ;
    RECT 8.83 87.195 16.37 89.015 ;
    LAYER Via34 ;
    RECT 8.83 121.125 16.37 121.905 ;
    LAYER Via34 ;
    RECT 8.83 126.185 16.37 126.965 ;
    LAYER Via34 ;
    RECT 8.83 131.245 16.37 132.025 ;
    LAYER Via34 ;
    RECT 8.83 136.305 16.37 137.085 ;
    LAYER Via34 ;
    RECT 8.83 141.365 16.37 142.145 ;
    LAYER Via34 ;
    RECT 8.83 146.425 16.37 147.205 ;
    LAYER Via34 ;
    RECT 8.83 149.875 16.37 150.655 ;
    END
  #BEGINEXT "VSI SIGNATURE 1.0"
    #CREATOR "Artisan Components, Inc." ;
    #DATE "2001-04-10" ;
    #REVISION "1.0" ;
    #ENDEXT
  END ram_128x16A

MACRO ram_256x16A
  CLASS RING ;
  FOREIGN ram_256x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 598.22 BY 189.235 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 309.98 17.2 311.08 18.3 ;
      LAYER Metal2 ;
      RECT 309.98 17.2 311.08 18.3 ;
      LAYER Metal3 ;
      RECT 309.98 17.2 311.08 18.3 ;
      LAYER Metal4 ;
      RECT 309.98 17.2 311.08 18.3 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 306.32 17.2 307.42 18.3 ;
      LAYER Metal2 ;
      RECT 306.32 17.2 307.42 18.3 ;
      LAYER Metal3 ;
      RECT 306.32 17.2 307.42 18.3 ;
      LAYER Metal4 ;
      RECT 306.32 17.2 307.42 18.3 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 301.18 17.2 302.28 18.3 ;
      LAYER Metal2 ;
      RECT 301.18 17.2 302.28 18.3 ;
      LAYER Metal3 ;
      RECT 301.18 17.2 302.28 18.3 ;
      LAYER Metal4 ;
      RECT 301.18 17.2 302.28 18.3 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 297.52 17.2 298.62 18.3 ;
      LAYER Metal2 ;
      RECT 297.52 17.2 298.62 18.3 ;
      LAYER Metal3 ;
      RECT 297.52 17.2 298.62 18.3 ;
      LAYER Metal4 ;
      RECT 297.52 17.2 298.62 18.3 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 288.72 17.2 289.82 18.3 ;
      LAYER Metal2 ;
      RECT 288.72 17.2 289.82 18.3 ;
      LAYER Metal3 ;
      RECT 288.72 17.2 289.82 18.3 ;
      LAYER Metal4 ;
      RECT 288.72 17.2 289.82 18.3 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 283.58 17.2 284.68 18.3 ;
      LAYER Metal2 ;
      RECT 283.58 17.2 284.68 18.3 ;
      LAYER Metal3 ;
      RECT 283.58 17.2 284.68 18.3 ;
      LAYER Metal4 ;
      RECT 283.58 17.2 284.68 18.3 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 279.92 17.2 281.02 18.3 ;
      LAYER Metal2 ;
      RECT 279.92 17.2 281.02 18.3 ;
      LAYER Metal3 ;
      RECT 279.92 17.2 281.02 18.3 ;
      LAYER Metal4 ;
      RECT 279.92 17.2 281.02 18.3 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 271.12 17.2 272.22 18.3 ;
      LAYER Metal2 ;
      RECT 271.12 17.2 272.22 18.3 ;
      LAYER Metal3 ;
      RECT 271.12 17.2 272.22 18.3 ;
      LAYER Metal4 ;
      RECT 271.12 17.2 272.22 18.3 ;
      END
    END A[7]
  PIN CEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 318.68 17.2 319.78 18.3 ;
      LAYER Metal2 ;
      RECT 318.68 17.2 319.78 18.3 ;
      LAYER Metal3 ;
      RECT 318.68 17.2 319.78 18.3 ;
      LAYER Metal4 ;
      RECT 318.68 17.2 319.78 18.3 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
      RECT 333.21 17.2 334.31 18.3 ;
      LAYER Metal2 ;
      RECT 333.21 17.2 334.31 18.3 ;
      LAYER Metal3 ;
      RECT 333.21 17.2 334.31 18.3 ;
      LAYER Metal4 ;
      RECT 333.21 17.2 334.31 18.3 ;
      END
    END CLK
  PIN D[0]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal2 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal3 ;
      RECT 45.46 17.2 46.56 18.3 ;
      LAYER Metal4 ;
      RECT 45.46 17.2 46.56 18.3 ;
      END
    END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 419.48 17.2 420.58 18.3 ;
      LAYER Metal2 ;
      RECT 419.48 17.2 420.58 18.3 ;
      LAYER Metal3 ;
      RECT 419.48 17.2 420.58 18.3 ;
      LAYER Metal4 ;
      RECT 419.48 17.2 420.58 18.3 ;
      END
    END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 430.3 17.2 431.4 18.3 ;
      LAYER Metal2 ;
      RECT 430.3 17.2 431.4 18.3 ;
      LAYER Metal3 ;
      RECT 430.3 17.2 431.4 18.3 ;
      LAYER Metal4 ;
      RECT 430.3 17.2 431.4 18.3 ;
      END
    END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 480.16 17.2 481.26 18.3 ;
      LAYER Metal2 ;
      RECT 480.16 17.2 481.26 18.3 ;
      LAYER Metal3 ;
      RECT 480.16 17.2 481.26 18.3 ;
      LAYER Metal4 ;
      RECT 480.16 17.2 481.26 18.3 ;
      END
    END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 490.98 17.2 492.08 18.3 ;
      LAYER Metal2 ;
      RECT 490.98 17.2 492.08 18.3 ;
      LAYER Metal3 ;
      RECT 490.98 17.2 492.08 18.3 ;
      LAYER Metal4 ;
      RECT 490.98 17.2 492.08 18.3 ;
      END
    END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 540.84 17.2 541.94 18.3 ;
      LAYER Metal2 ;
      RECT 540.84 17.2 541.94 18.3 ;
      LAYER Metal3 ;
      RECT 540.84 17.2 541.94 18.3 ;
      LAYER Metal4 ;
      RECT 540.84 17.2 541.94 18.3 ;
      END
    END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 551.66 17.2 552.76 18.3 ;
      LAYER Metal2 ;
      RECT 551.66 17.2 552.76 18.3 ;
      LAYER Metal3 ;
      RECT 551.66 17.2 552.76 18.3 ;
      LAYER Metal4 ;
      RECT 551.66 17.2 552.76 18.3 ;
      END
    END D[15]
  PIN D[1]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal2 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal3 ;
      RECT 56.28 17.2 57.38 18.3 ;
      LAYER Metal4 ;
      RECT 56.28 17.2 57.38 18.3 ;
      END
    END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal2 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal3 ;
      RECT 106.14 17.2 107.24 18.3 ;
      LAYER Metal4 ;
      RECT 106.14 17.2 107.24 18.3 ;
      END
    END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal2 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal3 ;
      RECT 116.96 17.2 118.06 18.3 ;
      LAYER Metal4 ;
      RECT 116.96 17.2 118.06 18.3 ;
      END
    END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal2 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal3 ;
      RECT 166.82 17.2 167.92 18.3 ;
      LAYER Metal4 ;
      RECT 166.82 17.2 167.92 18.3 ;
      END
    END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal2 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal3 ;
      RECT 177.64 17.2 178.74 18.3 ;
      LAYER Metal4 ;
      RECT 177.64 17.2 178.74 18.3 ;
      END
    END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal2 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal3 ;
      RECT 227.5 17.2 228.6 18.3 ;
      LAYER Metal4 ;
      RECT 227.5 17.2 228.6 18.3 ;
      END
    END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal2 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal3 ;
      RECT 238.32 17.2 239.42 18.3 ;
      LAYER Metal4 ;
      RECT 238.32 17.2 239.42 18.3 ;
      END
    END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 358.8 17.2 359.9 18.3 ;
      LAYER Metal2 ;
      RECT 358.8 17.2 359.9 18.3 ;
      LAYER Metal3 ;
      RECT 358.8 17.2 359.9 18.3 ;
      LAYER Metal4 ;
      RECT 358.8 17.2 359.9 18.3 ;
      END
    END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 369.62 17.2 370.72 18.3 ;
      LAYER Metal2 ;
      RECT 369.62 17.2 370.72 18.3 ;
      LAYER Metal3 ;
      RECT 369.62 17.2 370.72 18.3 ;
      LAYER Metal4 ;
      RECT 369.62 17.2 370.72 18.3 ;
      END
    END D[9]
  PIN OEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 330.2 17.2 331.3 18.3 ;
      LAYER Metal2 ;
      RECT 330.2 17.2 331.3 18.3 ;
      LAYER Metal3 ;
      RECT 330.2 17.2 331.3 18.3 ;
      LAYER Metal4 ;
      RECT 330.2 17.2 331.3 18.3 ;
      END
    END OEN
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal2 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal3 ;
      RECT 39.98 17.2 41.08 18.3 ;
      LAYER Metal4 ;
      RECT 39.98 17.2 41.08 18.3 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 414.2 17.2 415.3 18.3 ;
      LAYER Metal2 ;
      RECT 414.2 17.2 415.3 18.3 ;
      LAYER Metal3 ;
      RECT 414.2 17.2 415.3 18.3 ;
      LAYER Metal4 ;
      RECT 414.2 17.2 415.3 18.3 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 435.58 17.2 436.68 18.3 ;
      LAYER Metal2 ;
      RECT 435.58 17.2 436.68 18.3 ;
      LAYER Metal3 ;
      RECT 435.58 17.2 436.68 18.3 ;
      LAYER Metal4 ;
      RECT 435.58 17.2 436.68 18.3 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 474.88 17.2 475.98 18.3 ;
      LAYER Metal2 ;
      RECT 474.88 17.2 475.98 18.3 ;
      LAYER Metal3 ;
      RECT 474.88 17.2 475.98 18.3 ;
      LAYER Metal4 ;
      RECT 474.88 17.2 475.98 18.3 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 496.26 17.2 497.36 18.3 ;
      LAYER Metal2 ;
      RECT 496.26 17.2 497.36 18.3 ;
      LAYER Metal3 ;
      RECT 496.26 17.2 497.36 18.3 ;
      LAYER Metal4 ;
      RECT 496.26 17.2 497.36 18.3 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 535.56 17.2 536.66 18.3 ;
      LAYER Metal2 ;
      RECT 535.56 17.2 536.66 18.3 ;
      LAYER Metal3 ;
      RECT 535.56 17.2 536.66 18.3 ;
      LAYER Metal4 ;
      RECT 535.56 17.2 536.66 18.3 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 557.04 17.2 558.14 18.3 ;
      LAYER Metal2 ;
      RECT 557.04 17.2 558.14 18.3 ;
      LAYER Metal3 ;
      RECT 557.04 17.2 558.14 18.3 ;
      LAYER Metal4 ;
      RECT 557.04 17.2 558.14 18.3 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal2 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal3 ;
      RECT 61.56 17.2 62.66 18.3 ;
      LAYER Metal4 ;
      RECT 61.56 17.2 62.66 18.3 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal2 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal3 ;
      RECT 100.86 17.2 101.96 18.3 ;
      LAYER Metal4 ;
      RECT 100.86 17.2 101.96 18.3 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal2 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal3 ;
      RECT 122.24 17.2 123.34 18.3 ;
      LAYER Metal4 ;
      RECT 122.24 17.2 123.34 18.3 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal2 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal3 ;
      RECT 161.54 17.2 162.64 18.3 ;
      LAYER Metal4 ;
      RECT 161.54 17.2 162.64 18.3 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal2 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal3 ;
      RECT 182.92 17.2 184.02 18.3 ;
      LAYER Metal4 ;
      RECT 182.92 17.2 184.02 18.3 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal2 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal3 ;
      RECT 222.22 17.2 223.32 18.3 ;
      LAYER Metal4 ;
      RECT 222.22 17.2 223.32 18.3 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal2 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal3 ;
      RECT 243.6 17.2 244.7 18.3 ;
      LAYER Metal4 ;
      RECT 243.6 17.2 244.7 18.3 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 353.52 17.2 354.62 18.3 ;
      LAYER Metal2 ;
      RECT 353.52 17.2 354.62 18.3 ;
      LAYER Metal3 ;
      RECT 353.52 17.2 354.62 18.3 ;
      LAYER Metal4 ;
      RECT 353.52 17.2 354.62 18.3 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 374.9 17.2 376 18.3 ;
      LAYER Metal2 ;
      RECT 374.9 17.2 376 18.3 ;
      LAYER Metal3 ;
      RECT 374.9 17.2 376 18.3 ;
      LAYER Metal4 ;
      RECT 374.9 17.2 376 18.3 ;
      END
    END Q[9]
  PIN WEN
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 321.56 17.2 322.66 18.3 ;
      LAYER Metal2 ;
      RECT 321.56 17.2 322.66 18.3 ;
      LAYER Metal3 ;
      RECT 321.56 17.2 322.66 18.3 ;
      LAYER Metal4 ;
      RECT 321.56 17.2 322.66 18.3 ;
      END
    END WEN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 598.22 181.235 0 189.235 ;
      LAYER Metal5 ;
      RECT 0 0 598.22 8 ;
      LAYER Metal3 ;
      RECT 598.22 181.235 0 189.235 ;
      LAYER Metal3 ;
      RECT 0 0 598.22 8 ;
      LAYER Metal4 ;
      RECT 590.22 0 598.22 189.235 ;
      LAYER Metal4 ;
      RECT 0 189.235 8 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 589.62 172.635 8.6 180.635 ;
      LAYER Metal5 ;
      RECT 8.6 8.6 589.62 16.6 ;
      LAYER Metal3 ;
      RECT 589.62 172.635 8.6 180.635 ;
      LAYER Metal3 ;
      RECT 8.6 8.6 589.62 16.6 ;
      LAYER Metal4 ;
      RECT 581.62 8.6 589.62 180.635 ;
      LAYER Metal4 ;
      RECT 8.6 180.635 16.6 8.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Metal1 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Metal2 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Metal3 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Metal4 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Via12 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Via23 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Via34 ;
    RECT 17.2 17.2 581.02 172.035 ;
    LAYER Via34 ;
    RECT 581.85 172.865 589.39 180.405 ;
    LAYER Via34 ;
    RECT 8.83 8.83 16.37 16.37 ;
    LAYER Via34 ;
    RECT 581.85 8.83 589.39 16.37 ;
    LAYER Via34 ;
    RECT 8.83 172.865 16.37 180.405 ;
    LAYER Via34 ;
    RECT 590.45 181.465 597.99 189.005 ;
    LAYER Via34 ;
    RECT 0.23 0.23 7.77 7.77 ;
    LAYER Via34 ;
    RECT 590.45 0.23 597.99 7.77 ;
    LAYER Via34 ;
    RECT 0.23 181.465 7.77 189.005 ;
    LAYER Metal4 ;
    RECT 18.62 172.035 19.7 189.235 ;
    LAYER Metal4 ;
    RECT 24.1 172.035 25.26 189.235 ;
    LAYER Metal4 ;
    RECT 26.06 172.035 27.22 189.235 ;
    LAYER Metal4 ;
    RECT 31.46 172.035 32.62 189.235 ;
    LAYER Metal4 ;
    RECT 33.42 172.035 34.58 189.235 ;
    LAYER Metal4 ;
    RECT 38.82 172.035 39.98 189.235 ;
    LAYER Metal4 ;
    RECT 40.78 172.035 41.94 189.235 ;
    LAYER Metal4 ;
    RECT 46.18 172.035 47.34 189.235 ;
    LAYER Metal4 ;
    RECT 48.14 172.035 49.3 189.235 ;
    LAYER Metal4 ;
    RECT 53.54 172.035 54.7 189.235 ;
    LAYER Metal4 ;
    RECT 55.5 172.035 56.66 189.235 ;
    LAYER Metal4 ;
    RECT 60.9 172.035 62.06 189.235 ;
    LAYER Metal4 ;
    RECT 62.86 172.035 64.02 189.235 ;
    LAYER Metal4 ;
    RECT 68.26 172.035 69.42 189.235 ;
    LAYER Metal4 ;
    RECT 70.22 172.035 71.38 189.235 ;
    LAYER Metal4 ;
    RECT 75.62 172.035 76.78 189.235 ;
    LAYER Metal4 ;
    RECT 77.58 172.035 78.74 189.235 ;
    LAYER Metal4 ;
    RECT 84.78 172.035 85.94 189.235 ;
    LAYER Metal4 ;
    RECT 86.74 172.035 87.9 189.235 ;
    LAYER Metal4 ;
    RECT 92.14 172.035 93.3 189.235 ;
    LAYER Metal4 ;
    RECT 94.1 172.035 95.26 189.235 ;
    LAYER Metal4 ;
    RECT 99.5 172.035 100.66 189.235 ;
    LAYER Metal4 ;
    RECT 101.46 172.035 102.62 189.235 ;
    LAYER Metal4 ;
    RECT 106.86 172.035 108.02 189.235 ;
    LAYER Metal4 ;
    RECT 108.82 172.035 109.98 189.235 ;
    LAYER Metal4 ;
    RECT 114.22 172.035 115.38 189.235 ;
    LAYER Metal4 ;
    RECT 116.18 172.035 117.34 189.235 ;
    LAYER Metal4 ;
    RECT 121.58 172.035 122.74 189.235 ;
    LAYER Metal4 ;
    RECT 123.54 172.035 124.7 189.235 ;
    LAYER Metal4 ;
    RECT 128.94 172.035 130.1 189.235 ;
    LAYER Metal4 ;
    RECT 130.9 172.035 132.06 189.235 ;
    LAYER Metal4 ;
    RECT 136.3 172.035 137.46 189.235 ;
    LAYER Metal4 ;
    RECT 138.26 172.035 139.42 189.235 ;
    LAYER Metal4 ;
    RECT 145.46 172.035 146.62 189.235 ;
    LAYER Metal4 ;
    RECT 147.42 172.035 148.58 189.235 ;
    LAYER Metal4 ;
    RECT 152.82 172.035 153.98 189.235 ;
    LAYER Metal4 ;
    RECT 154.78 172.035 155.94 189.235 ;
    LAYER Metal4 ;
    RECT 160.18 172.035 161.34 189.235 ;
    LAYER Metal4 ;
    RECT 162.14 172.035 163.3 189.235 ;
    LAYER Metal4 ;
    RECT 167.54 172.035 168.7 189.235 ;
    LAYER Metal4 ;
    RECT 169.5 172.035 170.66 189.235 ;
    LAYER Metal4 ;
    RECT 174.9 172.035 176.06 189.235 ;
    LAYER Metal4 ;
    RECT 176.86 172.035 178.02 189.235 ;
    LAYER Metal4 ;
    RECT 182.26 172.035 183.42 189.235 ;
    LAYER Metal4 ;
    RECT 184.22 172.035 185.38 189.235 ;
    LAYER Metal4 ;
    RECT 189.62 172.035 190.78 189.235 ;
    LAYER Metal4 ;
    RECT 191.58 172.035 192.74 189.235 ;
    LAYER Metal4 ;
    RECT 196.98 172.035 198.14 189.235 ;
    LAYER Metal4 ;
    RECT 198.94 172.035 200.1 189.235 ;
    LAYER Metal4 ;
    RECT 206.14 172.035 207.3 189.235 ;
    LAYER Metal4 ;
    RECT 208.1 172.035 209.26 189.235 ;
    LAYER Metal4 ;
    RECT 213.5 172.035 214.66 189.235 ;
    LAYER Metal4 ;
    RECT 215.46 172.035 216.62 189.235 ;
    LAYER Metal4 ;
    RECT 220.86 172.035 222.02 189.235 ;
    LAYER Metal4 ;
    RECT 222.82 172.035 223.98 189.235 ;
    LAYER Metal4 ;
    RECT 228.22 172.035 229.38 189.235 ;
    LAYER Metal4 ;
    RECT 230.18 172.035 231.34 189.235 ;
    LAYER Metal4 ;
    RECT 235.58 172.035 236.74 189.235 ;
    LAYER Metal4 ;
    RECT 237.54 172.035 238.7 189.235 ;
    LAYER Metal4 ;
    RECT 242.94 172.035 244.1 189.235 ;
    LAYER Metal4 ;
    RECT 244.9 172.035 246.06 189.235 ;
    LAYER Metal4 ;
    RECT 250.3 172.035 251.46 189.235 ;
    LAYER Metal4 ;
    RECT 252.26 172.035 253.42 189.235 ;
    LAYER Metal4 ;
    RECT 257.66 172.035 258.82 189.235 ;
    LAYER Metal4 ;
    RECT 259.62 172.035 260.78 189.235 ;
    LAYER Metal4 ;
    RECT 264.96 172.035 266.64 189.235 ;
    LAYER Metal4 ;
    RECT 269.36 172.035 271.04 189.235 ;
    LAYER Metal4 ;
    RECT 273.76 172.035 275.44 189.235 ;
    LAYER Metal4 ;
    RECT 278.16 172.035 279.84 189.235 ;
    LAYER Metal4 ;
    RECT 282.56 172.035 284.24 189.235 ;
    LAYER Metal4 ;
    RECT 286.96 172.035 288.64 189.235 ;
    LAYER Metal4 ;
    RECT 291.36 172.035 293.04 189.235 ;
    LAYER Metal4 ;
    RECT 295.76 172.035 297.44 189.235 ;
    LAYER Metal4 ;
    RECT 300.16 172.035 301.84 189.235 ;
    LAYER Metal4 ;
    RECT 304.56 172.035 306.24 189.235 ;
    LAYER Metal4 ;
    RECT 308.96 172.035 310.64 189.235 ;
    LAYER Metal4 ;
    RECT 314.72 172.035 315.92 189.235 ;
    LAYER Metal4 ;
    RECT 319.66 172.035 321.68 189.235 ;
    LAYER Metal4 ;
    RECT 325.42 172.035 327.44 189.235 ;
    LAYER Metal4 ;
    RECT 330.12 172.035 331.4 189.235 ;
    LAYER Metal4 ;
    RECT 333.7 172.035 335.14 189.235 ;
    LAYER Metal4 ;
    RECT 337.44 172.035 338.6 189.235 ;
    LAYER Metal4 ;
    RECT 339.4 172.035 340.56 189.235 ;
    LAYER Metal4 ;
    RECT 344.8 172.035 345.96 189.235 ;
    LAYER Metal4 ;
    RECT 346.76 172.035 347.92 189.235 ;
    LAYER Metal4 ;
    RECT 352.16 172.035 353.32 189.235 ;
    LAYER Metal4 ;
    RECT 354.12 172.035 355.28 189.235 ;
    LAYER Metal4 ;
    RECT 359.52 172.035 360.68 189.235 ;
    LAYER Metal4 ;
    RECT 361.48 172.035 362.64 189.235 ;
    LAYER Metal4 ;
    RECT 366.88 172.035 368.04 189.235 ;
    LAYER Metal4 ;
    RECT 368.84 172.035 370 189.235 ;
    LAYER Metal4 ;
    RECT 374.24 172.035 375.4 189.235 ;
    LAYER Metal4 ;
    RECT 376.2 172.035 377.36 189.235 ;
    LAYER Metal4 ;
    RECT 381.6 172.035 382.76 189.235 ;
    LAYER Metal4 ;
    RECT 383.56 172.035 384.72 189.235 ;
    LAYER Metal4 ;
    RECT 388.96 172.035 390.12 189.235 ;
    LAYER Metal4 ;
    RECT 390.92 172.035 392.08 189.235 ;
    LAYER Metal4 ;
    RECT 398.12 172.035 399.28 189.235 ;
    LAYER Metal4 ;
    RECT 400.08 172.035 401.24 189.235 ;
    LAYER Metal4 ;
    RECT 405.48 172.035 406.64 189.235 ;
    LAYER Metal4 ;
    RECT 407.44 172.035 408.6 189.235 ;
    LAYER Metal4 ;
    RECT 412.84 172.035 414 189.235 ;
    LAYER Metal4 ;
    RECT 414.8 172.035 415.96 189.235 ;
    LAYER Metal4 ;
    RECT 420.2 172.035 421.36 189.235 ;
    LAYER Metal4 ;
    RECT 422.16 172.035 423.32 189.235 ;
    LAYER Metal4 ;
    RECT 427.56 172.035 428.72 189.235 ;
    LAYER Metal4 ;
    RECT 429.52 172.035 430.68 189.235 ;
    LAYER Metal4 ;
    RECT 434.92 172.035 436.08 189.235 ;
    LAYER Metal4 ;
    RECT 436.88 172.035 438.04 189.235 ;
    LAYER Metal4 ;
    RECT 442.28 172.035 443.44 189.235 ;
    LAYER Metal4 ;
    RECT 444.24 172.035 445.4 189.235 ;
    LAYER Metal4 ;
    RECT 449.64 172.035 450.8 189.235 ;
    LAYER Metal4 ;
    RECT 451.6 172.035 452.76 189.235 ;
    LAYER Metal4 ;
    RECT 458.8 172.035 459.96 189.235 ;
    LAYER Metal4 ;
    RECT 460.76 172.035 461.92 189.235 ;
    LAYER Metal4 ;
    RECT 466.16 172.035 467.32 189.235 ;
    LAYER Metal4 ;
    RECT 468.12 172.035 469.28 189.235 ;
    LAYER Metal4 ;
    RECT 473.52 172.035 474.68 189.235 ;
    LAYER Metal4 ;
    RECT 475.48 172.035 476.64 189.235 ;
    LAYER Metal4 ;
    RECT 480.88 172.035 482.04 189.235 ;
    LAYER Metal4 ;
    RECT 482.84 172.035 484 189.235 ;
    LAYER Metal4 ;
    RECT 488.24 172.035 489.4 189.235 ;
    LAYER Metal4 ;
    RECT 490.2 172.035 491.36 189.235 ;
    LAYER Metal4 ;
    RECT 495.6 172.035 496.76 189.235 ;
    LAYER Metal4 ;
    RECT 497.56 172.035 498.72 189.235 ;
    LAYER Metal4 ;
    RECT 502.96 172.035 504.12 189.235 ;
    LAYER Metal4 ;
    RECT 504.92 172.035 506.08 189.235 ;
    LAYER Metal4 ;
    RECT 510.32 172.035 511.48 189.235 ;
    LAYER Metal4 ;
    RECT 512.28 172.035 513.44 189.235 ;
    LAYER Metal4 ;
    RECT 519.48 172.035 520.64 189.235 ;
    LAYER Metal4 ;
    RECT 521.44 172.035 522.6 189.235 ;
    LAYER Metal4 ;
    RECT 526.84 172.035 528 189.235 ;
    LAYER Metal4 ;
    RECT 528.8 172.035 529.96 189.235 ;
    LAYER Metal4 ;
    RECT 534.2 172.035 535.36 189.235 ;
    LAYER Metal4 ;
    RECT 536.16 172.035 537.32 189.235 ;
    LAYER Metal4 ;
    RECT 541.56 172.035 542.72 189.235 ;
    LAYER Metal4 ;
    RECT 543.52 172.035 544.68 189.235 ;
    LAYER Metal4 ;
    RECT 548.92 172.035 550.08 189.235 ;
    LAYER Metal4 ;
    RECT 550.88 172.035 552.04 189.235 ;
    LAYER Metal4 ;
    RECT 556.28 172.035 557.44 189.235 ;
    LAYER Metal4 ;
    RECT 558.24 172.035 559.4 189.235 ;
    LAYER Metal4 ;
    RECT 563.64 172.035 564.8 189.235 ;
    LAYER Metal4 ;
    RECT 565.6 172.035 566.76 189.235 ;
    LAYER Metal4 ;
    RECT 571 172.035 572.16 189.235 ;
    LAYER Metal4 ;
    RECT 572.96 172.035 574.12 189.235 ;
    LAYER Metal4 ;
    RECT 578.52 172.035 579.6 189.235 ;
    LAYER Metal4 ;
    RECT 18.02 17.2 19.12 0 ;
    LAYER Metal4 ;
    RECT 24.1 17.2 27.22 0 ;
    LAYER Metal4 ;
    RECT 31.46 17.2 34.58 0 ;
    LAYER Metal4 ;
    RECT 38.18 17.2 39.52 0 ;
    LAYER Metal4 ;
    RECT 47.02 17.2 49.4 0 ;
    LAYER Metal4 ;
    RECT 53.44 17.2 55.82 0 ;
    LAYER Metal4 ;
    RECT 63.32 17.2 64.66 0 ;
    LAYER Metal4 ;
    RECT 68.26 17.2 71.38 0 ;
    LAYER Metal4 ;
    RECT 75.62 17.2 78.74 0 ;
    LAYER Metal4 ;
    RECT 84.78 17.2 87.9 0 ;
    LAYER Metal4 ;
    RECT 92.14 17.2 95.26 0 ;
    LAYER Metal4 ;
    RECT 98.86 17.2 100.2 0 ;
    LAYER Metal4 ;
    RECT 107.7 17.2 110.08 0 ;
    LAYER Metal4 ;
    RECT 114.12 17.2 116.5 0 ;
    LAYER Metal4 ;
    RECT 124 17.2 125.34 0 ;
    LAYER Metal4 ;
    RECT 128.94 17.2 132.06 0 ;
    LAYER Metal4 ;
    RECT 136.3 17.2 139.42 0 ;
    LAYER Metal4 ;
    RECT 145.46 17.2 148.58 0 ;
    LAYER Metal4 ;
    RECT 152.82 17.2 155.94 0 ;
    LAYER Metal4 ;
    RECT 159.54 17.2 160.88 0 ;
    LAYER Metal4 ;
    RECT 168.38 17.2 170.76 0 ;
    LAYER Metal4 ;
    RECT 174.8 17.2 177.18 0 ;
    LAYER Metal4 ;
    RECT 184.68 17.2 186.02 0 ;
    LAYER Metal4 ;
    RECT 189.62 17.2 192.74 0 ;
    LAYER Metal4 ;
    RECT 196.98 17.2 200.1 0 ;
    LAYER Metal4 ;
    RECT 206.14 17.2 209.26 0 ;
    LAYER Metal4 ;
    RECT 213.5 17.2 216.62 0 ;
    LAYER Metal4 ;
    RECT 220.22 17.2 221.56 0 ;
    LAYER Metal4 ;
    RECT 229.06 17.2 231.44 0 ;
    LAYER Metal4 ;
    RECT 235.48 17.2 237.86 0 ;
    LAYER Metal4 ;
    RECT 245.36 17.2 246.7 0 ;
    LAYER Metal4 ;
    RECT 250.3 17.2 253.42 0 ;
    LAYER Metal4 ;
    RECT 257.66 17.2 260.78 0 ;
    LAYER Metal4 ;
    RECT 268.28 17.2 269.92 0 ;
    LAYER Metal4 ;
    RECT 274.98 17.2 278.78 0 ;
    LAYER Metal4 ;
    RECT 285.88 17.2 287.52 0 ;
    LAYER Metal4 ;
    RECT 292.58 17.2 296.38 0 ;
    LAYER Metal4 ;
    RECT 303.48 17.2 305.12 0 ;
    LAYER Metal4 ;
    RECT 312.83 17.2 313.37 0 ;
    LAYER Metal4 ;
    RECT 314.41 17.2 315.41 0 ;
    LAYER Metal4 ;
    RECT 320.24 17.2 321.1 0 ;
    LAYER Metal4 ;
    RECT 326 17.2 326.86 0 ;
    LAYER Metal4 ;
    RECT 337.44 17.2 340.56 0 ;
    LAYER Metal4 ;
    RECT 344.8 17.2 347.92 0 ;
    LAYER Metal4 ;
    RECT 351.52 17.2 352.86 0 ;
    LAYER Metal4 ;
    RECT 360.36 17.2 362.74 0 ;
    LAYER Metal4 ;
    RECT 366.78 17.2 369.16 0 ;
    LAYER Metal4 ;
    RECT 376.66 17.2 378 0 ;
    LAYER Metal4 ;
    RECT 381.6 17.2 384.72 0 ;
    LAYER Metal4 ;
    RECT 388.96 17.2 392.08 0 ;
    LAYER Metal4 ;
    RECT 398.12 17.2 401.24 0 ;
    LAYER Metal4 ;
    RECT 405.48 17.2 408.6 0 ;
    LAYER Metal4 ;
    RECT 412.2 17.2 413.54 0 ;
    LAYER Metal4 ;
    RECT 421.04 17.2 423.42 0 ;
    LAYER Metal4 ;
    RECT 427.46 17.2 429.84 0 ;
    LAYER Metal4 ;
    RECT 437.34 17.2 438.68 0 ;
    LAYER Metal4 ;
    RECT 442.28 17.2 445.4 0 ;
    LAYER Metal4 ;
    RECT 449.64 17.2 452.76 0 ;
    LAYER Metal4 ;
    RECT 458.8 17.2 461.92 0 ;
    LAYER Metal4 ;
    RECT 466.16 17.2 469.28 0 ;
    LAYER Metal4 ;
    RECT 472.88 17.2 474.22 0 ;
    LAYER Metal4 ;
    RECT 481.72 17.2 484.1 0 ;
    LAYER Metal4 ;
    RECT 488.14 17.2 490.52 0 ;
    LAYER Metal4 ;
    RECT 498.02 17.2 499.36 0 ;
    LAYER Metal4 ;
    RECT 502.96 17.2 506.08 0 ;
    LAYER Metal4 ;
    RECT 510.32 17.2 513.44 0 ;
    LAYER Metal4 ;
    RECT 519.48 17.2 522.6 0 ;
    LAYER Metal4 ;
    RECT 526.84 17.2 529.96 0 ;
    LAYER Metal4 ;
    RECT 533.56 17.2 534.9 0 ;
    LAYER Metal4 ;
    RECT 542.4 17.2 544.78 0 ;
    LAYER Metal4 ;
    RECT 548.82 17.2 551.2 0 ;
    LAYER Metal4 ;
    RECT 558.7 17.2 560.04 0 ;
    LAYER Metal4 ;
    RECT 563.64 17.2 566.76 0 ;
    LAYER Metal4 ;
    RECT 571 17.2 574.12 0 ;
    LAYER Metal4 ;
    RECT 579.1 17.2 580.2 0 ;
    LAYER Metal3 ;
    RECT 581.02 22.22 598.22 23.22 ;
    LAYER Metal3 ;
    RECT 581.02 35.14 598.22 36.04 ;
    LAYER Metal3 ;
    RECT 581.02 48.245 598.22 48.845 ;
    LAYER Metal3 ;
    RECT 581.02 52.605 598.22 53.505 ;
    LAYER Metal3 ;
    RECT 581.02 73.205 598.22 73.805 ;
    LAYER Metal3 ;
    RECT 581.02 82.685 598.22 84.285 ;
    LAYER Metal3 ;
    RECT 581.02 90.11 598.22 94.61 ;
    LAYER Metal3 ;
    RECT 581.02 95.21 598.22 103.61 ;
    LAYER Metal3 ;
    RECT 581.02 105.875 598.22 109.575 ;
    LAYER Metal3 ;
    RECT 581.02 110.19 598.22 114.19 ;
    LAYER Metal3 ;
    RECT 581.02 123.595 598.22 124.495 ;
    LAYER Metal3 ;
    RECT 581.02 128.655 598.22 129.555 ;
    LAYER Metal3 ;
    RECT 581.02 133.715 598.22 134.615 ;
    LAYER Metal3 ;
    RECT 581.02 138.775 598.22 139.675 ;
    LAYER Metal3 ;
    RECT 581.02 143.835 598.22 144.735 ;
    LAYER Metal3 ;
    RECT 581.02 148.895 598.22 149.795 ;
    LAYER Metal3 ;
    RECT 581.02 153.955 598.22 154.855 ;
    LAYER Metal3 ;
    RECT 581.02 159.015 598.22 159.915 ;
    LAYER Metal3 ;
    RECT 581.02 164.345 598.22 165.245 ;
    LAYER Metal3 ;
    RECT 581.02 168.245 598.22 169.145 ;
    LAYER Metal3 ;
    RECT 17.2 22.22 0 23.22 ;
    LAYER Metal3 ;
    RECT 17.2 35.14 0 36.04 ;
    LAYER Metal3 ;
    RECT 17.2 48.245 0 48.845 ;
    LAYER Metal3 ;
    RECT 17.2 52.605 0 53.505 ;
    LAYER Metal3 ;
    RECT 17.2 73.205 0 73.805 ;
    LAYER Metal3 ;
    RECT 17.2 82.685 0 84.285 ;
    LAYER Metal3 ;
    RECT 17.2 90.11 0 94.61 ;
    LAYER Metal3 ;
    RECT 17.2 95.21 0 103.61 ;
    LAYER Metal3 ;
    RECT 17.2 105.875 0 109.575 ;
    LAYER Metal3 ;
    RECT 17.2 110.19 0 114.19 ;
    LAYER Metal3 ;
    RECT 17.2 123.595 0 124.495 ;
    LAYER Metal3 ;
    RECT 17.2 128.655 0 129.555 ;
    LAYER Metal3 ;
    RECT 17.2 133.715 0 134.615 ;
    LAYER Metal3 ;
    RECT 17.2 138.775 0 139.675 ;
    LAYER Metal3 ;
    RECT 17.2 143.835 0 144.735 ;
    LAYER Metal3 ;
    RECT 17.2 148.895 0 149.795 ;
    LAYER Metal3 ;
    RECT 17.2 153.955 0 154.855 ;
    LAYER Metal3 ;
    RECT 17.2 159.015 0 159.915 ;
    LAYER Metal3 ;
    RECT 17.2 164.345 0 165.245 ;
    LAYER Metal3 ;
    RECT 17.2 168.245 0 169.145 ;
    LAYER Metal4 ;
    RECT 20.42 172.035 21.7 180.635 ;
    LAYER Metal4 ;
    RECT 22.38 172.035 23.54 180.635 ;
    LAYER Metal4 ;
    RECT 27.78 172.035 28.94 180.635 ;
    LAYER Metal4 ;
    RECT 29.74 172.035 30.9 180.635 ;
    LAYER Metal4 ;
    RECT 35.14 172.035 36.3 180.635 ;
    LAYER Metal4 ;
    RECT 37.1 172.035 38.26 180.635 ;
    LAYER Metal4 ;
    RECT 42.5 172.035 43.66 180.635 ;
    LAYER Metal4 ;
    RECT 44.46 172.035 45.62 180.635 ;
    LAYER Metal4 ;
    RECT 49.86 172.035 51.02 180.635 ;
    LAYER Metal4 ;
    RECT 51.82 172.035 52.98 180.635 ;
    LAYER Metal4 ;
    RECT 57.22 172.035 58.38 180.635 ;
    LAYER Metal4 ;
    RECT 59.18 172.035 60.34 180.635 ;
    LAYER Metal4 ;
    RECT 64.58 172.035 65.74 180.635 ;
    LAYER Metal4 ;
    RECT 66.54 172.035 67.7 180.635 ;
    LAYER Metal4 ;
    RECT 71.94 172.035 73.1 180.635 ;
    LAYER Metal4 ;
    RECT 73.9 172.035 75.06 180.635 ;
    LAYER Metal4 ;
    RECT 79.3 172.035 80.46 180.635 ;
    LAYER Metal4 ;
    RECT 81.21 172.035 82.31 180.635 ;
    LAYER Metal4 ;
    RECT 83.06 172.035 84.22 180.635 ;
    LAYER Metal4 ;
    RECT 88.46 172.035 89.62 180.635 ;
    LAYER Metal4 ;
    RECT 90.42 172.035 91.58 180.635 ;
    LAYER Metal4 ;
    RECT 95.82 172.035 96.98 180.635 ;
    LAYER Metal4 ;
    RECT 97.78 172.035 98.94 180.635 ;
    LAYER Metal4 ;
    RECT 103.18 172.035 104.34 180.635 ;
    LAYER Metal4 ;
    RECT 105.14 172.035 106.3 180.635 ;
    LAYER Metal4 ;
    RECT 110.54 172.035 111.7 180.635 ;
    LAYER Metal4 ;
    RECT 112.5 172.035 113.66 180.635 ;
    LAYER Metal4 ;
    RECT 117.9 172.035 119.06 180.635 ;
    LAYER Metal4 ;
    RECT 119.86 172.035 121.02 180.635 ;
    LAYER Metal4 ;
    RECT 125.26 172.035 126.42 180.635 ;
    LAYER Metal4 ;
    RECT 127.22 172.035 128.38 180.635 ;
    LAYER Metal4 ;
    RECT 132.62 172.035 133.78 180.635 ;
    LAYER Metal4 ;
    RECT 134.58 172.035 135.74 180.635 ;
    LAYER Metal4 ;
    RECT 139.98 172.035 141.14 180.635 ;
    LAYER Metal4 ;
    RECT 141.89 172.035 142.99 180.635 ;
    LAYER Metal4 ;
    RECT 143.74 172.035 144.9 180.635 ;
    LAYER Metal4 ;
    RECT 149.14 172.035 150.3 180.635 ;
    LAYER Metal4 ;
    RECT 151.1 172.035 152.26 180.635 ;
    LAYER Metal4 ;
    RECT 156.5 172.035 157.66 180.635 ;
    LAYER Metal4 ;
    RECT 158.46 172.035 159.62 180.635 ;
    LAYER Metal4 ;
    RECT 163.86 172.035 165.02 180.635 ;
    LAYER Metal4 ;
    RECT 165.82 172.035 166.98 180.635 ;
    LAYER Metal4 ;
    RECT 171.22 172.035 172.38 180.635 ;
    LAYER Metal4 ;
    RECT 173.18 172.035 174.34 180.635 ;
    LAYER Metal4 ;
    RECT 178.58 172.035 179.74 180.635 ;
    LAYER Metal4 ;
    RECT 180.54 172.035 181.7 180.635 ;
    LAYER Metal4 ;
    RECT 185.94 172.035 187.1 180.635 ;
    LAYER Metal4 ;
    RECT 187.9 172.035 189.06 180.635 ;
    LAYER Metal4 ;
    RECT 193.3 172.035 194.46 180.635 ;
    LAYER Metal4 ;
    RECT 195.26 172.035 196.42 180.635 ;
    LAYER Metal4 ;
    RECT 200.66 172.035 201.82 180.635 ;
    LAYER Metal4 ;
    RECT 202.57 172.035 203.67 180.635 ;
    LAYER Metal4 ;
    RECT 204.42 172.035 205.58 180.635 ;
    LAYER Metal4 ;
    RECT 209.82 172.035 210.98 180.635 ;
    LAYER Metal4 ;
    RECT 211.78 172.035 212.94 180.635 ;
    LAYER Metal4 ;
    RECT 217.18 172.035 218.34 180.635 ;
    LAYER Metal4 ;
    RECT 219.14 172.035 220.3 180.635 ;
    LAYER Metal4 ;
    RECT 224.54 172.035 225.7 180.635 ;
    LAYER Metal4 ;
    RECT 226.5 172.035 227.66 180.635 ;
    LAYER Metal4 ;
    RECT 231.9 172.035 233.06 180.635 ;
    LAYER Metal4 ;
    RECT 233.86 172.035 235.02 180.635 ;
    LAYER Metal4 ;
    RECT 239.26 172.035 240.42 180.635 ;
    LAYER Metal4 ;
    RECT 241.22 172.035 242.38 180.635 ;
    LAYER Metal4 ;
    RECT 246.62 172.035 247.78 180.635 ;
    LAYER Metal4 ;
    RECT 248.58 172.035 249.74 180.635 ;
    LAYER Metal4 ;
    RECT 253.98 172.035 255.14 180.635 ;
    LAYER Metal4 ;
    RECT 255.94 172.035 257.1 180.635 ;
    LAYER Metal4 ;
    RECT 261.34 172.035 262.5 180.635 ;
    LAYER Metal4 ;
    RECT 263.25 172.035 264.35 180.635 ;
    LAYER Metal4 ;
    RECT 267.1 172.035 268.9 180.635 ;
    LAYER Metal4 ;
    RECT 271.56 172.035 273.24 180.635 ;
    LAYER Metal4 ;
    RECT 275.96 172.035 277.64 180.635 ;
    LAYER Metal4 ;
    RECT 280.36 172.035 282.04 180.635 ;
    LAYER Metal4 ;
    RECT 284.76 172.035 286.44 180.635 ;
    LAYER Metal4 ;
    RECT 289.16 172.035 290.84 180.635 ;
    LAYER Metal4 ;
    RECT 293.56 172.035 295.24 180.635 ;
    LAYER Metal4 ;
    RECT 297.96 172.035 299.64 180.635 ;
    LAYER Metal4 ;
    RECT 302.36 172.035 304.04 180.635 ;
    LAYER Metal4 ;
    RECT 306.76 172.035 308.44 180.635 ;
    LAYER Metal4 ;
    RECT 311.1 172.035 314.1 180.635 ;
    LAYER Metal4 ;
    RECT 316.78 172.035 318.8 180.635 ;
    LAYER Metal4 ;
    RECT 322.54 172.035 324.56 180.635 ;
    LAYER Metal4 ;
    RECT 328.3 172.035 329.5 180.635 ;
    LAYER Metal4 ;
    RECT 331.96 172.035 333.24 180.635 ;
    LAYER Metal4 ;
    RECT 335.72 172.035 336.88 180.635 ;
    LAYER Metal4 ;
    RECT 341.12 172.035 342.28 180.635 ;
    LAYER Metal4 ;
    RECT 343.08 172.035 344.24 180.635 ;
    LAYER Metal4 ;
    RECT 348.48 172.035 349.64 180.635 ;
    LAYER Metal4 ;
    RECT 350.44 172.035 351.6 180.635 ;
    LAYER Metal4 ;
    RECT 355.84 172.035 357 180.635 ;
    LAYER Metal4 ;
    RECT 357.8 172.035 358.96 180.635 ;
    LAYER Metal4 ;
    RECT 363.2 172.035 364.36 180.635 ;
    LAYER Metal4 ;
    RECT 365.16 172.035 366.32 180.635 ;
    LAYER Metal4 ;
    RECT 370.56 172.035 371.72 180.635 ;
    LAYER Metal4 ;
    RECT 372.52 172.035 373.68 180.635 ;
    LAYER Metal4 ;
    RECT 377.92 172.035 379.08 180.635 ;
    LAYER Metal4 ;
    RECT 379.88 172.035 381.04 180.635 ;
    LAYER Metal4 ;
    RECT 385.28 172.035 386.44 180.635 ;
    LAYER Metal4 ;
    RECT 387.24 172.035 388.4 180.635 ;
    LAYER Metal4 ;
    RECT 392.64 172.035 393.8 180.635 ;
    LAYER Metal4 ;
    RECT 394.55 172.035 395.65 180.635 ;
    LAYER Metal4 ;
    RECT 396.4 172.035 397.56 180.635 ;
    LAYER Metal4 ;
    RECT 401.8 172.035 402.96 180.635 ;
    LAYER Metal4 ;
    RECT 403.76 172.035 404.92 180.635 ;
    LAYER Metal4 ;
    RECT 409.16 172.035 410.32 180.635 ;
    LAYER Metal4 ;
    RECT 411.12 172.035 412.28 180.635 ;
    LAYER Metal4 ;
    RECT 416.52 172.035 417.68 180.635 ;
    LAYER Metal4 ;
    RECT 418.48 172.035 419.64 180.635 ;
    LAYER Metal4 ;
    RECT 423.88 172.035 425.04 180.635 ;
    LAYER Metal4 ;
    RECT 425.84 172.035 427 180.635 ;
    LAYER Metal4 ;
    RECT 431.24 172.035 432.4 180.635 ;
    LAYER Metal4 ;
    RECT 433.2 172.035 434.36 180.635 ;
    LAYER Metal4 ;
    RECT 438.6 172.035 439.76 180.635 ;
    LAYER Metal4 ;
    RECT 440.56 172.035 441.72 180.635 ;
    LAYER Metal4 ;
    RECT 445.96 172.035 447.12 180.635 ;
    LAYER Metal4 ;
    RECT 447.92 172.035 449.08 180.635 ;
    LAYER Metal4 ;
    RECT 453.32 172.035 454.48 180.635 ;
    LAYER Metal4 ;
    RECT 455.23 172.035 456.33 180.635 ;
    LAYER Metal4 ;
    RECT 457.08 172.035 458.24 180.635 ;
    LAYER Metal4 ;
    RECT 462.48 172.035 463.64 180.635 ;
    LAYER Metal4 ;
    RECT 464.44 172.035 465.6 180.635 ;
    LAYER Metal4 ;
    RECT 469.84 172.035 471 180.635 ;
    LAYER Metal4 ;
    RECT 471.8 172.035 472.96 180.635 ;
    LAYER Metal4 ;
    RECT 477.2 172.035 478.36 180.635 ;
    LAYER Metal4 ;
    RECT 479.16 172.035 480.32 180.635 ;
    LAYER Metal4 ;
    RECT 484.56 172.035 485.72 180.635 ;
    LAYER Metal4 ;
    RECT 486.52 172.035 487.68 180.635 ;
    LAYER Metal4 ;
    RECT 491.92 172.035 493.08 180.635 ;
    LAYER Metal4 ;
    RECT 493.88 172.035 495.04 180.635 ;
    LAYER Metal4 ;
    RECT 499.28 172.035 500.44 180.635 ;
    LAYER Metal4 ;
    RECT 501.24 172.035 502.4 180.635 ;
    LAYER Metal4 ;
    RECT 506.64 172.035 507.8 180.635 ;
    LAYER Metal4 ;
    RECT 508.6 172.035 509.76 180.635 ;
    LAYER Metal4 ;
    RECT 514 172.035 515.16 180.635 ;
    LAYER Metal4 ;
    RECT 515.91 172.035 517.01 180.635 ;
    LAYER Metal4 ;
    RECT 517.76 172.035 518.92 180.635 ;
    LAYER Metal4 ;
    RECT 523.16 172.035 524.32 180.635 ;
    LAYER Metal4 ;
    RECT 525.12 172.035 526.28 180.635 ;
    LAYER Metal4 ;
    RECT 530.52 172.035 531.68 180.635 ;
    LAYER Metal4 ;
    RECT 532.48 172.035 533.64 180.635 ;
    LAYER Metal4 ;
    RECT 537.88 172.035 539.04 180.635 ;
    LAYER Metal4 ;
    RECT 539.84 172.035 541 180.635 ;
    LAYER Metal4 ;
    RECT 545.24 172.035 546.4 180.635 ;
    LAYER Metal4 ;
    RECT 547.2 172.035 548.36 180.635 ;
    LAYER Metal4 ;
    RECT 552.6 172.035 553.76 180.635 ;
    LAYER Metal4 ;
    RECT 554.56 172.035 555.72 180.635 ;
    LAYER Metal4 ;
    RECT 559.96 172.035 561.12 180.635 ;
    LAYER Metal4 ;
    RECT 561.92 172.035 563.08 180.635 ;
    LAYER Metal4 ;
    RECT 567.32 172.035 568.48 180.635 ;
    LAYER Metal4 ;
    RECT 569.28 172.035 570.44 180.635 ;
    LAYER Metal4 ;
    RECT 574.68 172.035 575.84 180.635 ;
    LAYER Metal4 ;
    RECT 576.52 172.035 577.8 180.635 ;
    LAYER Metal4 ;
    RECT 19.58 17.2 20.78 8.6 ;
    LAYER Metal4 ;
    RECT 21.48 17.2 22.48 8.6 ;
    LAYER Metal4 ;
    RECT 27.78 17.2 30.9 8.6 ;
    LAYER Metal4 ;
    RECT 36.2 17.2 37.2 8.6 ;
    LAYER Metal4 ;
    RECT 43.1 17.2 44.32 8.6 ;
    LAYER Metal4 ;
    RECT 50.82 17.2 52.02 8.6 ;
    LAYER Metal4 ;
    RECT 58.52 17.2 59.74 8.6 ;
    LAYER Metal4 ;
    RECT 65.64 17.2 66.64 8.6 ;
    LAYER Metal4 ;
    RECT 71.94 17.2 75.06 8.6 ;
    LAYER Metal4 ;
    RECT 80.36 17.2 81.36 8.6 ;
    LAYER Metal4 ;
    RECT 82.16 17.2 83.16 8.6 ;
    LAYER Metal4 ;
    RECT 88.46 17.2 91.58 8.6 ;
    LAYER Metal4 ;
    RECT 96.88 17.2 97.88 8.6 ;
    LAYER Metal4 ;
    RECT 103.78 17.2 105 8.6 ;
    LAYER Metal4 ;
    RECT 111.5 17.2 112.7 8.6 ;
    LAYER Metal4 ;
    RECT 119.2 17.2 120.42 8.6 ;
    LAYER Metal4 ;
    RECT 126.32 17.2 127.32 8.6 ;
    LAYER Metal4 ;
    RECT 132.62 17.2 135.74 8.6 ;
    LAYER Metal4 ;
    RECT 141.04 17.2 142.04 8.6 ;
    LAYER Metal4 ;
    RECT 142.84 17.2 143.84 8.6 ;
    LAYER Metal4 ;
    RECT 149.14 17.2 152.26 8.6 ;
    LAYER Metal4 ;
    RECT 157.56 17.2 158.56 8.6 ;
    LAYER Metal4 ;
    RECT 164.46 17.2 165.68 8.6 ;
    LAYER Metal4 ;
    RECT 172.18 17.2 173.38 8.6 ;
    LAYER Metal4 ;
    RECT 179.88 17.2 181.1 8.6 ;
    LAYER Metal4 ;
    RECT 187 17.2 188 8.6 ;
    LAYER Metal4 ;
    RECT 193.3 17.2 196.42 8.6 ;
    LAYER Metal4 ;
    RECT 201.72 17.2 202.72 8.6 ;
    LAYER Metal4 ;
    RECT 203.52 17.2 204.52 8.6 ;
    LAYER Metal4 ;
    RECT 209.82 17.2 212.94 8.6 ;
    LAYER Metal4 ;
    RECT 218.24 17.2 219.24 8.6 ;
    LAYER Metal4 ;
    RECT 225.14 17.2 226.36 8.6 ;
    LAYER Metal4 ;
    RECT 232.86 17.2 234.06 8.6 ;
    LAYER Metal4 ;
    RECT 240.56 17.2 241.78 8.6 ;
    LAYER Metal4 ;
    RECT 247.68 17.2 248.68 8.6 ;
    LAYER Metal4 ;
    RECT 253.98 17.2 257.1 8.6 ;
    LAYER Metal4 ;
    RECT 262.4 17.2 263.4 8.6 ;
    LAYER Metal4 ;
    RECT 264.2 17.2 265.2 8.6 ;
    LAYER Metal4 ;
    RECT 265.91 17.2 267.51 8.6 ;
    LAYER Metal4 ;
    RECT 272.68 17.2 274.32 8.6 ;
    LAYER Metal4 ;
    RECT 281.48 17.2 283.12 8.6 ;
    LAYER Metal4 ;
    RECT 290.28 17.2 291.92 8.6 ;
    LAYER Metal4 ;
    RECT 299.08 17.2 300.72 8.6 ;
    LAYER Metal4 ;
    RECT 307.88 17.2 309.52 8.6 ;
    LAYER Metal4 ;
    RECT 317.36 17.2 318.22 8.6 ;
    LAYER Metal4 ;
    RECT 323.12 17.2 323.98 8.6 ;
    LAYER Metal4 ;
    RECT 328.88 17.2 329.74 8.6 ;
    LAYER Metal4 ;
    RECT 331.77 17.2 332.75 8.6 ;
    LAYER Metal4 ;
    RECT 334.82 17.2 335.82 8.6 ;
    LAYER Metal4 ;
    RECT 341.12 17.2 344.24 8.6 ;
    LAYER Metal4 ;
    RECT 349.54 17.2 350.54 8.6 ;
    LAYER Metal4 ;
    RECT 356.44 17.2 357.66 8.6 ;
    LAYER Metal4 ;
    RECT 364.16 17.2 365.36 8.6 ;
    LAYER Metal4 ;
    RECT 371.86 17.2 373.08 8.6 ;
    LAYER Metal4 ;
    RECT 378.98 17.2 379.98 8.6 ;
    LAYER Metal4 ;
    RECT 385.28 17.2 388.4 8.6 ;
    LAYER Metal4 ;
    RECT 393.7 17.2 394.7 8.6 ;
    LAYER Metal4 ;
    RECT 395.5 17.2 396.5 8.6 ;
    LAYER Metal4 ;
    RECT 401.8 17.2 404.92 8.6 ;
    LAYER Metal4 ;
    RECT 410.22 17.2 411.22 8.6 ;
    LAYER Metal4 ;
    RECT 417.12 17.2 418.34 8.6 ;
    LAYER Metal4 ;
    RECT 424.84 17.2 426.04 8.6 ;
    LAYER Metal4 ;
    RECT 432.54 17.2 433.76 8.6 ;
    LAYER Metal4 ;
    RECT 439.66 17.2 440.66 8.6 ;
    LAYER Metal4 ;
    RECT 445.96 17.2 449.08 8.6 ;
    LAYER Metal4 ;
    RECT 454.38 17.2 455.38 8.6 ;
    LAYER Metal4 ;
    RECT 456.18 17.2 457.18 8.6 ;
    LAYER Metal4 ;
    RECT 462.48 17.2 465.6 8.6 ;
    LAYER Metal4 ;
    RECT 470.9 17.2 471.9 8.6 ;
    LAYER Metal4 ;
    RECT 477.8 17.2 479.02 8.6 ;
    LAYER Metal4 ;
    RECT 485.52 17.2 486.72 8.6 ;
    LAYER Metal4 ;
    RECT 493.22 17.2 494.44 8.6 ;
    LAYER Metal4 ;
    RECT 500.34 17.2 501.34 8.6 ;
    LAYER Metal4 ;
    RECT 506.64 17.2 509.76 8.6 ;
    LAYER Metal4 ;
    RECT 515.06 17.2 516.06 8.6 ;
    LAYER Metal4 ;
    RECT 516.86 17.2 517.86 8.6 ;
    LAYER Metal4 ;
    RECT 523.16 17.2 526.28 8.6 ;
    LAYER Metal4 ;
    RECT 531.58 17.2 532.58 8.6 ;
    LAYER Metal4 ;
    RECT 538.48 17.2 539.7 8.6 ;
    LAYER Metal4 ;
    RECT 546.2 17.2 547.4 8.6 ;
    LAYER Metal4 ;
    RECT 553.9 17.2 555.12 8.6 ;
    LAYER Metal4 ;
    RECT 561.02 17.2 562.02 8.6 ;
    LAYER Metal4 ;
    RECT 567.32 17.2 570.44 8.6 ;
    LAYER Metal4 ;
    RECT 575.74 17.2 576.74 8.6 ;
    LAYER Metal4 ;
    RECT 577.44 17.2 578.64 8.6 ;
    LAYER Metal3 ;
    RECT 581.02 28.715 589.62 30.115 ;
    LAYER Metal3 ;
    RECT 581.02 54.775 589.62 57.275 ;
    LAYER Metal3 ;
    RECT 581.02 63.17 589.62 67.97 ;
    LAYER Metal3 ;
    RECT 581.02 74.265 589.62 74.865 ;
    LAYER Metal3 ;
    RECT 581.02 87.105 589.62 89.105 ;
    LAYER Metal3 ;
    RECT 581.02 121.065 589.62 121.965 ;
    LAYER Metal3 ;
    RECT 581.02 126.125 589.62 127.025 ;
    LAYER Metal3 ;
    RECT 581.02 131.185 589.62 132.085 ;
    LAYER Metal3 ;
    RECT 581.02 136.245 589.62 137.145 ;
    LAYER Metal3 ;
    RECT 581.02 141.305 589.62 142.205 ;
    LAYER Metal3 ;
    RECT 581.02 146.365 589.62 147.265 ;
    LAYER Metal3 ;
    RECT 581.02 151.425 589.62 152.325 ;
    LAYER Metal3 ;
    RECT 581.02 156.485 589.62 157.385 ;
    LAYER Metal3 ;
    RECT 581.02 161.545 589.62 162.445 ;
    LAYER Metal3 ;
    RECT 581.02 166.605 589.62 167.505 ;
    LAYER Metal3 ;
    RECT 581.02 170.055 589.62 170.955 ;
    LAYER Metal3 ;
    RECT 17.2 28.715 8.6 30.115 ;
    LAYER Metal3 ;
    RECT 17.2 54.775 8.6 57.275 ;
    LAYER Metal3 ;
    RECT 17.2 63.17 8.6 67.97 ;
    LAYER Metal3 ;
    RECT 17.2 74.265 8.6 74.865 ;
    LAYER Metal3 ;
    RECT 17.2 87.105 8.6 89.105 ;
    LAYER Metal3 ;
    RECT 17.2 121.065 8.6 121.965 ;
    LAYER Metal3 ;
    RECT 17.2 126.125 8.6 127.025 ;
    LAYER Metal3 ;
    RECT 17.2 131.185 8.6 132.085 ;
    LAYER Metal3 ;
    RECT 17.2 136.245 8.6 137.145 ;
    LAYER Metal3 ;
    RECT 17.2 141.305 8.6 142.205 ;
    LAYER Metal3 ;
    RECT 17.2 146.365 8.6 147.265 ;
    LAYER Metal3 ;
    RECT 17.2 151.425 8.6 152.325 ;
    LAYER Metal3 ;
    RECT 17.2 156.485 8.6 157.385 ;
    LAYER Metal3 ;
    RECT 17.2 161.545 8.6 162.445 ;
    LAYER Metal3 ;
    RECT 17.2 166.605 8.6 167.505 ;
    LAYER Metal3 ;
    RECT 17.2 170.055 8.6 170.955 ;
    LAYER Via34 ;
    RECT 18.77 181.465 19.55 189.005 ;
    LAYER Via34 ;
    RECT 24.29 181.465 25.07 189.005 ;
    LAYER Via34 ;
    RECT 26.25 181.465 27.03 189.005 ;
    LAYER Via34 ;
    RECT 31.65 181.465 32.43 189.005 ;
    LAYER Via34 ;
    RECT 33.61 181.465 34.39 189.005 ;
    LAYER Via34 ;
    RECT 39.01 181.465 39.79 189.005 ;
    LAYER Via34 ;
    RECT 40.97 181.465 41.75 189.005 ;
    LAYER Via34 ;
    RECT 46.37 181.465 47.15 189.005 ;
    LAYER Via34 ;
    RECT 48.33 181.465 49.11 189.005 ;
    LAYER Via34 ;
    RECT 53.73 181.465 54.51 189.005 ;
    LAYER Via34 ;
    RECT 55.69 181.465 56.47 189.005 ;
    LAYER Via34 ;
    RECT 61.09 181.465 61.87 189.005 ;
    LAYER Via34 ;
    RECT 63.05 181.465 63.83 189.005 ;
    LAYER Via34 ;
    RECT 68.45 181.465 69.23 189.005 ;
    LAYER Via34 ;
    RECT 70.41 181.465 71.19 189.005 ;
    LAYER Via34 ;
    RECT 75.81 181.465 76.59 189.005 ;
    LAYER Via34 ;
    RECT 77.77 181.465 78.55 189.005 ;
    LAYER Via34 ;
    RECT 84.97 181.465 85.75 189.005 ;
    LAYER Via34 ;
    RECT 86.93 181.465 87.71 189.005 ;
    LAYER Via34 ;
    RECT 92.33 181.465 93.11 189.005 ;
    LAYER Via34 ;
    RECT 94.29 181.465 95.07 189.005 ;
    LAYER Via34 ;
    RECT 99.69 181.465 100.47 189.005 ;
    LAYER Via34 ;
    RECT 101.65 181.465 102.43 189.005 ;
    LAYER Via34 ;
    RECT 107.05 181.465 107.83 189.005 ;
    LAYER Via34 ;
    RECT 109.01 181.465 109.79 189.005 ;
    LAYER Via34 ;
    RECT 114.41 181.465 115.19 189.005 ;
    LAYER Via34 ;
    RECT 116.37 181.465 117.15 189.005 ;
    LAYER Via34 ;
    RECT 121.77 181.465 122.55 189.005 ;
    LAYER Via34 ;
    RECT 123.73 181.465 124.51 189.005 ;
    LAYER Via34 ;
    RECT 129.13 181.465 129.91 189.005 ;
    LAYER Via34 ;
    RECT 131.09 181.465 131.87 189.005 ;
    LAYER Via34 ;
    RECT 136.49 181.465 137.27 189.005 ;
    LAYER Via34 ;
    RECT 138.45 181.465 139.23 189.005 ;
    LAYER Via34 ;
    RECT 145.65 181.465 146.43 189.005 ;
    LAYER Via34 ;
    RECT 147.61 181.465 148.39 189.005 ;
    LAYER Via34 ;
    RECT 153.01 181.465 153.79 189.005 ;
    LAYER Via34 ;
    RECT 154.97 181.465 155.75 189.005 ;
    LAYER Via34 ;
    RECT 160.37 181.465 161.15 189.005 ;
    LAYER Via34 ;
    RECT 162.33 181.465 163.11 189.005 ;
    LAYER Via34 ;
    RECT 167.73 181.465 168.51 189.005 ;
    LAYER Via34 ;
    RECT 169.69 181.465 170.47 189.005 ;
    LAYER Via34 ;
    RECT 175.09 181.465 175.87 189.005 ;
    LAYER Via34 ;
    RECT 177.05 181.465 177.83 189.005 ;
    LAYER Via34 ;
    RECT 182.45 181.465 183.23 189.005 ;
    LAYER Via34 ;
    RECT 184.41 181.465 185.19 189.005 ;
    LAYER Via34 ;
    RECT 189.81 181.465 190.59 189.005 ;
    LAYER Via34 ;
    RECT 191.77 181.465 192.55 189.005 ;
    LAYER Via34 ;
    RECT 197.17 181.465 197.95 189.005 ;
    LAYER Via34 ;
    RECT 199.13 181.465 199.91 189.005 ;
    LAYER Via34 ;
    RECT 206.33 181.465 207.11 189.005 ;
    LAYER Via34 ;
    RECT 208.29 181.465 209.07 189.005 ;
    LAYER Via34 ;
    RECT 213.69 181.465 214.47 189.005 ;
    LAYER Via34 ;
    RECT 215.65 181.465 216.43 189.005 ;
    LAYER Via34 ;
    RECT 221.05 181.465 221.83 189.005 ;
    LAYER Via34 ;
    RECT 223.01 181.465 223.79 189.005 ;
    LAYER Via34 ;
    RECT 228.41 181.465 229.19 189.005 ;
    LAYER Via34 ;
    RECT 230.37 181.465 231.15 189.005 ;
    LAYER Via34 ;
    RECT 235.77 181.465 236.55 189.005 ;
    LAYER Via34 ;
    RECT 237.73 181.465 238.51 189.005 ;
    LAYER Via34 ;
    RECT 243.13 181.465 243.91 189.005 ;
    LAYER Via34 ;
    RECT 245.09 181.465 245.87 189.005 ;
    LAYER Via34 ;
    RECT 250.49 181.465 251.27 189.005 ;
    LAYER Via34 ;
    RECT 252.45 181.465 253.23 189.005 ;
    LAYER Via34 ;
    RECT 257.85 181.465 258.63 189.005 ;
    LAYER Via34 ;
    RECT 259.81 181.465 260.59 189.005 ;
    LAYER Via34 ;
    RECT 265.15 181.465 266.45 189.005 ;
    LAYER Via34 ;
    RECT 269.55 181.465 270.85 189.005 ;
    LAYER Via34 ;
    RECT 273.95 181.465 275.25 189.005 ;
    LAYER Via34 ;
    RECT 278.35 181.465 279.65 189.005 ;
    LAYER Via34 ;
    RECT 282.75 181.465 284.05 189.005 ;
    LAYER Via34 ;
    RECT 287.15 181.465 288.45 189.005 ;
    LAYER Via34 ;
    RECT 291.55 181.465 292.85 189.005 ;
    LAYER Via34 ;
    RECT 295.95 181.465 297.25 189.005 ;
    LAYER Via34 ;
    RECT 300.35 181.465 301.65 189.005 ;
    LAYER Via34 ;
    RECT 304.75 181.465 306.05 189.005 ;
    LAYER Via34 ;
    RECT 309.15 181.465 310.45 189.005 ;
    LAYER Via34 ;
    RECT 314.93 181.465 315.71 189.005 ;
    LAYER Via34 ;
    RECT 319.76 181.465 321.58 189.005 ;
    LAYER Via34 ;
    RECT 325.52 181.465 327.34 189.005 ;
    LAYER Via34 ;
    RECT 330.37 181.465 331.15 189.005 ;
    LAYER Via34 ;
    RECT 333.77 181.465 335.07 189.005 ;
    LAYER Via34 ;
    RECT 337.63 181.465 338.41 189.005 ;
    LAYER Via34 ;
    RECT 339.59 181.465 340.37 189.005 ;
    LAYER Via34 ;
    RECT 344.99 181.465 345.77 189.005 ;
    LAYER Via34 ;
    RECT 346.95 181.465 347.73 189.005 ;
    LAYER Via34 ;
    RECT 352.35 181.465 353.13 189.005 ;
    LAYER Via34 ;
    RECT 354.31 181.465 355.09 189.005 ;
    LAYER Via34 ;
    RECT 359.71 181.465 360.49 189.005 ;
    LAYER Via34 ;
    RECT 361.67 181.465 362.45 189.005 ;
    LAYER Via34 ;
    RECT 367.07 181.465 367.85 189.005 ;
    LAYER Via34 ;
    RECT 369.03 181.465 369.81 189.005 ;
    LAYER Via34 ;
    RECT 374.43 181.465 375.21 189.005 ;
    LAYER Via34 ;
    RECT 376.39 181.465 377.17 189.005 ;
    LAYER Via34 ;
    RECT 381.79 181.465 382.57 189.005 ;
    LAYER Via34 ;
    RECT 383.75 181.465 384.53 189.005 ;
    LAYER Via34 ;
    RECT 389.15 181.465 389.93 189.005 ;
    LAYER Via34 ;
    RECT 391.11 181.465 391.89 189.005 ;
    LAYER Via34 ;
    RECT 398.31 181.465 399.09 189.005 ;
    LAYER Via34 ;
    RECT 400.27 181.465 401.05 189.005 ;
    LAYER Via34 ;
    RECT 405.67 181.465 406.45 189.005 ;
    LAYER Via34 ;
    RECT 407.63 181.465 408.41 189.005 ;
    LAYER Via34 ;
    RECT 413.03 181.465 413.81 189.005 ;
    LAYER Via34 ;
    RECT 414.99 181.465 415.77 189.005 ;
    LAYER Via34 ;
    RECT 420.39 181.465 421.17 189.005 ;
    LAYER Via34 ;
    RECT 422.35 181.465 423.13 189.005 ;
    LAYER Via34 ;
    RECT 427.75 181.465 428.53 189.005 ;
    LAYER Via34 ;
    RECT 429.71 181.465 430.49 189.005 ;
    LAYER Via34 ;
    RECT 435.11 181.465 435.89 189.005 ;
    LAYER Via34 ;
    RECT 437.07 181.465 437.85 189.005 ;
    LAYER Via34 ;
    RECT 442.47 181.465 443.25 189.005 ;
    LAYER Via34 ;
    RECT 444.43 181.465 445.21 189.005 ;
    LAYER Via34 ;
    RECT 449.83 181.465 450.61 189.005 ;
    LAYER Via34 ;
    RECT 451.79 181.465 452.57 189.005 ;
    LAYER Via34 ;
    RECT 458.99 181.465 459.77 189.005 ;
    LAYER Via34 ;
    RECT 460.95 181.465 461.73 189.005 ;
    LAYER Via34 ;
    RECT 466.35 181.465 467.13 189.005 ;
    LAYER Via34 ;
    RECT 468.31 181.465 469.09 189.005 ;
    LAYER Via34 ;
    RECT 473.71 181.465 474.49 189.005 ;
    LAYER Via34 ;
    RECT 475.67 181.465 476.45 189.005 ;
    LAYER Via34 ;
    RECT 481.07 181.465 481.85 189.005 ;
    LAYER Via34 ;
    RECT 483.03 181.465 483.81 189.005 ;
    LAYER Via34 ;
    RECT 488.43 181.465 489.21 189.005 ;
    LAYER Via34 ;
    RECT 490.39 181.465 491.17 189.005 ;
    LAYER Via34 ;
    RECT 495.79 181.465 496.57 189.005 ;
    LAYER Via34 ;
    RECT 497.75 181.465 498.53 189.005 ;
    LAYER Via34 ;
    RECT 503.15 181.465 503.93 189.005 ;
    LAYER Via34 ;
    RECT 505.11 181.465 505.89 189.005 ;
    LAYER Via34 ;
    RECT 510.51 181.465 511.29 189.005 ;
    LAYER Via34 ;
    RECT 512.47 181.465 513.25 189.005 ;
    LAYER Via34 ;
    RECT 519.67 181.465 520.45 189.005 ;
    LAYER Via34 ;
    RECT 521.63 181.465 522.41 189.005 ;
    LAYER Via34 ;
    RECT 527.03 181.465 527.81 189.005 ;
    LAYER Via34 ;
    RECT 528.99 181.465 529.77 189.005 ;
    LAYER Via34 ;
    RECT 534.39 181.465 535.17 189.005 ;
    LAYER Via34 ;
    RECT 536.35 181.465 537.13 189.005 ;
    LAYER Via34 ;
    RECT 541.75 181.465 542.53 189.005 ;
    LAYER Via34 ;
    RECT 543.71 181.465 544.49 189.005 ;
    LAYER Via34 ;
    RECT 549.11 181.465 549.89 189.005 ;
    LAYER Via34 ;
    RECT 551.07 181.465 551.85 189.005 ;
    LAYER Via34 ;
    RECT 556.47 181.465 557.25 189.005 ;
    LAYER Via34 ;
    RECT 558.43 181.465 559.21 189.005 ;
    LAYER Via34 ;
    RECT 563.83 181.465 564.61 189.005 ;
    LAYER Via34 ;
    RECT 565.79 181.465 566.57 189.005 ;
    LAYER Via34 ;
    RECT 571.19 181.465 571.97 189.005 ;
    LAYER Via34 ;
    RECT 573.15 181.465 573.93 189.005 ;
    LAYER Via34 ;
    RECT 578.67 181.465 579.45 189.005 ;
    LAYER Via34 ;
    RECT 18.18 0.23 18.96 7.77 ;
    LAYER Via34 ;
    RECT 24.23 0.23 27.09 7.77 ;
    LAYER Via34 ;
    RECT 31.59 0.23 34.45 7.77 ;
    LAYER Via34 ;
    RECT 38.46 0.23 39.24 7.77 ;
    LAYER Via34 ;
    RECT 47.3 0.23 49.12 7.77 ;
    LAYER Via34 ;
    RECT 53.72 0.23 55.54 7.77 ;
    LAYER Via34 ;
    RECT 63.6 0.23 64.38 7.77 ;
    LAYER Via34 ;
    RECT 68.39 0.23 71.25 7.77 ;
    LAYER Via34 ;
    RECT 75.75 0.23 78.61 7.77 ;
    LAYER Via34 ;
    RECT 84.91 0.23 87.77 7.77 ;
    LAYER Via34 ;
    RECT 92.27 0.23 95.13 7.77 ;
    LAYER Via34 ;
    RECT 99.14 0.23 99.92 7.77 ;
    LAYER Via34 ;
    RECT 107.98 0.23 109.8 7.77 ;
    LAYER Via34 ;
    RECT 114.4 0.23 116.22 7.77 ;
    LAYER Via34 ;
    RECT 124.28 0.23 125.06 7.77 ;
    LAYER Via34 ;
    RECT 129.07 0.23 131.93 7.77 ;
    LAYER Via34 ;
    RECT 136.43 0.23 139.29 7.77 ;
    LAYER Via34 ;
    RECT 145.59 0.23 148.45 7.77 ;
    LAYER Via34 ;
    RECT 152.95 0.23 155.81 7.77 ;
    LAYER Via34 ;
    RECT 159.82 0.23 160.6 7.77 ;
    LAYER Via34 ;
    RECT 168.66 0.23 170.48 7.77 ;
    LAYER Via34 ;
    RECT 175.08 0.23 176.9 7.77 ;
    LAYER Via34 ;
    RECT 184.96 0.23 185.74 7.77 ;
    LAYER Via34 ;
    RECT 189.75 0.23 192.61 7.77 ;
    LAYER Via34 ;
    RECT 197.11 0.23 199.97 7.77 ;
    LAYER Via34 ;
    RECT 206.27 0.23 209.13 7.77 ;
    LAYER Via34 ;
    RECT 213.63 0.23 216.49 7.77 ;
    LAYER Via34 ;
    RECT 220.5 0.23 221.28 7.77 ;
    LAYER Via34 ;
    RECT 229.34 0.23 231.16 7.77 ;
    LAYER Via34 ;
    RECT 235.76 0.23 237.58 7.77 ;
    LAYER Via34 ;
    RECT 245.64 0.23 246.42 7.77 ;
    LAYER Via34 ;
    RECT 250.43 0.23 253.29 7.77 ;
    LAYER Via34 ;
    RECT 257.79 0.23 260.65 7.77 ;
    LAYER Via34 ;
    RECT 268.45 0.23 269.75 7.77 ;
    LAYER Via34 ;
    RECT 275.19 0.23 278.57 7.77 ;
    LAYER Via34 ;
    RECT 286.05 0.23 287.35 7.77 ;
    LAYER Via34 ;
    RECT 292.79 0.23 296.17 7.77 ;
    LAYER Via34 ;
    RECT 303.65 0.23 304.95 7.77 ;
    LAYER Via34 ;
    RECT 312.97 0.23 313.23 7.77 ;
    LAYER Via34 ;
    RECT 314.52 0.23 315.3 7.77 ;
    LAYER Via34 ;
    RECT 320.54 0.23 320.8 7.77 ;
    LAYER Via34 ;
    RECT 326.3 0.23 326.56 7.77 ;
    LAYER Via34 ;
    RECT 337.57 0.23 340.43 7.77 ;
    LAYER Via34 ;
    RECT 344.93 0.23 347.79 7.77 ;
    LAYER Via34 ;
    RECT 351.8 0.23 352.58 7.77 ;
    LAYER Via34 ;
    RECT 360.64 0.23 362.46 7.77 ;
    LAYER Via34 ;
    RECT 367.06 0.23 368.88 7.77 ;
    LAYER Via34 ;
    RECT 376.94 0.23 377.72 7.77 ;
    LAYER Via34 ;
    RECT 381.73 0.23 384.59 7.77 ;
    LAYER Via34 ;
    RECT 389.09 0.23 391.95 7.77 ;
    LAYER Via34 ;
    RECT 398.25 0.23 401.11 7.77 ;
    LAYER Via34 ;
    RECT 405.61 0.23 408.47 7.77 ;
    LAYER Via34 ;
    RECT 412.48 0.23 413.26 7.77 ;
    LAYER Via34 ;
    RECT 421.32 0.23 423.14 7.77 ;
    LAYER Via34 ;
    RECT 427.74 0.23 429.56 7.77 ;
    LAYER Via34 ;
    RECT 437.62 0.23 438.4 7.77 ;
    LAYER Via34 ;
    RECT 442.41 0.23 445.27 7.77 ;
    LAYER Via34 ;
    RECT 449.77 0.23 452.63 7.77 ;
    LAYER Via34 ;
    RECT 458.93 0.23 461.79 7.77 ;
    LAYER Via34 ;
    RECT 466.29 0.23 469.15 7.77 ;
    LAYER Via34 ;
    RECT 473.16 0.23 473.94 7.77 ;
    LAYER Via34 ;
    RECT 482 0.23 483.82 7.77 ;
    LAYER Via34 ;
    RECT 488.42 0.23 490.24 7.77 ;
    LAYER Via34 ;
    RECT 498.3 0.23 499.08 7.77 ;
    LAYER Via34 ;
    RECT 503.09 0.23 505.95 7.77 ;
    LAYER Via34 ;
    RECT 510.45 0.23 513.31 7.77 ;
    LAYER Via34 ;
    RECT 519.61 0.23 522.47 7.77 ;
    LAYER Via34 ;
    RECT 526.97 0.23 529.83 7.77 ;
    LAYER Via34 ;
    RECT 533.84 0.23 534.62 7.77 ;
    LAYER Via34 ;
    RECT 542.68 0.23 544.5 7.77 ;
    LAYER Via34 ;
    RECT 549.1 0.23 550.92 7.77 ;
    LAYER Via34 ;
    RECT 558.98 0.23 559.76 7.77 ;
    LAYER Via34 ;
    RECT 563.77 0.23 566.63 7.77 ;
    LAYER Via34 ;
    RECT 571.13 0.23 573.99 7.77 ;
    LAYER Via34 ;
    RECT 579.26 0.23 580.04 7.77 ;
    LAYER Via34 ;
    RECT 590.45 22.33 597.99 23.11 ;
    LAYER Via34 ;
    RECT 590.45 35.2 597.99 35.98 ;
    LAYER Via34 ;
    RECT 590.45 48.415 597.99 48.675 ;
    LAYER Via34 ;
    RECT 590.45 52.665 597.99 53.445 ;
    LAYER Via34 ;
    RECT 590.45 73.375 597.99 73.635 ;
    LAYER Via34 ;
    RECT 590.45 82.835 597.99 84.135 ;
    LAYER Via34 ;
    RECT 590.45 90.41 597.99 94.31 ;
    LAYER Via34 ;
    RECT 590.45 95.38 597.99 103.44 ;
    LAYER Via34 ;
    RECT 590.45 106.035 597.99 109.415 ;
    LAYER Via34 ;
    RECT 590.45 110.5 597.99 113.88 ;
    LAYER Via34 ;
    RECT 590.45 123.655 597.99 124.435 ;
    LAYER Via34 ;
    RECT 590.45 128.715 597.99 129.495 ;
    LAYER Via34 ;
    RECT 590.45 133.775 597.99 134.555 ;
    LAYER Via34 ;
    RECT 590.45 138.835 597.99 139.615 ;
    LAYER Via34 ;
    RECT 590.45 143.895 597.99 144.675 ;
    LAYER Via34 ;
    RECT 590.45 148.955 597.99 149.735 ;
    LAYER Via34 ;
    RECT 590.45 154.015 597.99 154.795 ;
    LAYER Via34 ;
    RECT 590.45 159.075 597.99 159.855 ;
    LAYER Via34 ;
    RECT 590.45 164.405 597.99 165.185 ;
    LAYER Via34 ;
    RECT 590.45 168.305 597.99 169.085 ;
    LAYER Via34 ;
    RECT 0.23 22.33 7.77 23.11 ;
    LAYER Via34 ;
    RECT 0.23 35.2 7.77 35.98 ;
    LAYER Via34 ;
    RECT 0.23 48.415 7.77 48.675 ;
    LAYER Via34 ;
    RECT 0.23 52.665 7.77 53.445 ;
    LAYER Via34 ;
    RECT 0.23 73.375 7.77 73.635 ;
    LAYER Via34 ;
    RECT 0.23 82.835 7.77 84.135 ;
    LAYER Via34 ;
    RECT 0.23 90.41 7.77 94.31 ;
    LAYER Via34 ;
    RECT 0.23 95.38 7.77 103.44 ;
    LAYER Via34 ;
    RECT 0.23 106.035 7.77 109.415 ;
    LAYER Via34 ;
    RECT 0.23 110.5 7.77 113.88 ;
    LAYER Via34 ;
    RECT 0.23 123.655 7.77 124.435 ;
    LAYER Via34 ;
    RECT 0.23 128.715 7.77 129.495 ;
    LAYER Via34 ;
    RECT 0.23 133.775 7.77 134.555 ;
    LAYER Via34 ;
    RECT 0.23 138.835 7.77 139.615 ;
    LAYER Via34 ;
    RECT 0.23 143.895 7.77 144.675 ;
    LAYER Via34 ;
    RECT 0.23 148.955 7.77 149.735 ;
    LAYER Via34 ;
    RECT 0.23 154.015 7.77 154.795 ;
    LAYER Via34 ;
    RECT 0.23 159.075 7.77 159.855 ;
    LAYER Via34 ;
    RECT 0.23 164.405 7.77 165.185 ;
    LAYER Via34 ;
    RECT 0.23 168.305 7.77 169.085 ;
    LAYER Via34 ;
    RECT 20.67 172.865 21.45 180.405 ;
    LAYER Via34 ;
    RECT 22.57 172.865 23.35 180.405 ;
    LAYER Via34 ;
    RECT 27.97 172.865 28.75 180.405 ;
    LAYER Via34 ;
    RECT 29.93 172.865 30.71 180.405 ;
    LAYER Via34 ;
    RECT 35.33 172.865 36.11 180.405 ;
    LAYER Via34 ;
    RECT 37.29 172.865 38.07 180.405 ;
    LAYER Via34 ;
    RECT 42.69 172.865 43.47 180.405 ;
    LAYER Via34 ;
    RECT 44.65 172.865 45.43 180.405 ;
    LAYER Via34 ;
    RECT 50.05 172.865 50.83 180.405 ;
    LAYER Via34 ;
    RECT 52.01 172.865 52.79 180.405 ;
    LAYER Via34 ;
    RECT 57.41 172.865 58.19 180.405 ;
    LAYER Via34 ;
    RECT 59.37 172.865 60.15 180.405 ;
    LAYER Via34 ;
    RECT 64.77 172.865 65.55 180.405 ;
    LAYER Via34 ;
    RECT 66.73 172.865 67.51 180.405 ;
    LAYER Via34 ;
    RECT 72.13 172.865 72.91 180.405 ;
    LAYER Via34 ;
    RECT 74.09 172.865 74.87 180.405 ;
    LAYER Via34 ;
    RECT 79.49 172.865 80.27 180.405 ;
    LAYER Via34 ;
    RECT 81.37 172.865 82.15 180.405 ;
    LAYER Via34 ;
    RECT 83.25 172.865 84.03 180.405 ;
    LAYER Via34 ;
    RECT 88.65 172.865 89.43 180.405 ;
    LAYER Via34 ;
    RECT 90.61 172.865 91.39 180.405 ;
    LAYER Via34 ;
    RECT 96.01 172.865 96.79 180.405 ;
    LAYER Via34 ;
    RECT 97.97 172.865 98.75 180.405 ;
    LAYER Via34 ;
    RECT 103.37 172.865 104.15 180.405 ;
    LAYER Via34 ;
    RECT 105.33 172.865 106.11 180.405 ;
    LAYER Via34 ;
    RECT 110.73 172.865 111.51 180.405 ;
    LAYER Via34 ;
    RECT 112.69 172.865 113.47 180.405 ;
    LAYER Via34 ;
    RECT 118.09 172.865 118.87 180.405 ;
    LAYER Via34 ;
    RECT 120.05 172.865 120.83 180.405 ;
    LAYER Via34 ;
    RECT 125.45 172.865 126.23 180.405 ;
    LAYER Via34 ;
    RECT 127.41 172.865 128.19 180.405 ;
    LAYER Via34 ;
    RECT 132.81 172.865 133.59 180.405 ;
    LAYER Via34 ;
    RECT 134.77 172.865 135.55 180.405 ;
    LAYER Via34 ;
    RECT 140.17 172.865 140.95 180.405 ;
    LAYER Via34 ;
    RECT 142.05 172.865 142.83 180.405 ;
    LAYER Via34 ;
    RECT 143.93 172.865 144.71 180.405 ;
    LAYER Via34 ;
    RECT 149.33 172.865 150.11 180.405 ;
    LAYER Via34 ;
    RECT 151.29 172.865 152.07 180.405 ;
    LAYER Via34 ;
    RECT 156.69 172.865 157.47 180.405 ;
    LAYER Via34 ;
    RECT 158.65 172.865 159.43 180.405 ;
    LAYER Via34 ;
    RECT 164.05 172.865 164.83 180.405 ;
    LAYER Via34 ;
    RECT 166.01 172.865 166.79 180.405 ;
    LAYER Via34 ;
    RECT 171.41 172.865 172.19 180.405 ;
    LAYER Via34 ;
    RECT 173.37 172.865 174.15 180.405 ;
    LAYER Via34 ;
    RECT 178.77 172.865 179.55 180.405 ;
    LAYER Via34 ;
    RECT 180.73 172.865 181.51 180.405 ;
    LAYER Via34 ;
    RECT 186.13 172.865 186.91 180.405 ;
    LAYER Via34 ;
    RECT 188.09 172.865 188.87 180.405 ;
    LAYER Via34 ;
    RECT 193.49 172.865 194.27 180.405 ;
    LAYER Via34 ;
    RECT 195.45 172.865 196.23 180.405 ;
    LAYER Via34 ;
    RECT 200.85 172.865 201.63 180.405 ;
    LAYER Via34 ;
    RECT 202.73 172.865 203.51 180.405 ;
    LAYER Via34 ;
    RECT 204.61 172.865 205.39 180.405 ;
    LAYER Via34 ;
    RECT 210.01 172.865 210.79 180.405 ;
    LAYER Via34 ;
    RECT 211.97 172.865 212.75 180.405 ;
    LAYER Via34 ;
    RECT 217.37 172.865 218.15 180.405 ;
    LAYER Via34 ;
    RECT 219.33 172.865 220.11 180.405 ;
    LAYER Via34 ;
    RECT 224.73 172.865 225.51 180.405 ;
    LAYER Via34 ;
    RECT 226.69 172.865 227.47 180.405 ;
    LAYER Via34 ;
    RECT 232.09 172.865 232.87 180.405 ;
    LAYER Via34 ;
    RECT 234.05 172.865 234.83 180.405 ;
    LAYER Via34 ;
    RECT 239.45 172.865 240.23 180.405 ;
    LAYER Via34 ;
    RECT 241.41 172.865 242.19 180.405 ;
    LAYER Via34 ;
    RECT 246.81 172.865 247.59 180.405 ;
    LAYER Via34 ;
    RECT 248.77 172.865 249.55 180.405 ;
    LAYER Via34 ;
    RECT 254.17 172.865 254.95 180.405 ;
    LAYER Via34 ;
    RECT 256.13 172.865 256.91 180.405 ;
    LAYER Via34 ;
    RECT 261.53 172.865 262.31 180.405 ;
    LAYER Via34 ;
    RECT 263.41 172.865 264.19 180.405 ;
    LAYER Via34 ;
    RECT 267.35 172.865 268.65 180.405 ;
    LAYER Via34 ;
    RECT 271.75 172.865 273.05 180.405 ;
    LAYER Via34 ;
    RECT 276.15 172.865 277.45 180.405 ;
    LAYER Via34 ;
    RECT 280.55 172.865 281.85 180.405 ;
    LAYER Via34 ;
    RECT 284.95 172.865 286.25 180.405 ;
    LAYER Via34 ;
    RECT 289.35 172.865 290.65 180.405 ;
    LAYER Via34 ;
    RECT 293.75 172.865 295.05 180.405 ;
    LAYER Via34 ;
    RECT 298.15 172.865 299.45 180.405 ;
    LAYER Via34 ;
    RECT 302.55 172.865 303.85 180.405 ;
    LAYER Via34 ;
    RECT 306.95 172.865 308.25 180.405 ;
    LAYER Via34 ;
    RECT 311.17 172.865 314.03 180.405 ;
    LAYER Via34 ;
    RECT 316.88 172.865 318.7 180.405 ;
    LAYER Via34 ;
    RECT 322.64 172.865 324.46 180.405 ;
    LAYER Via34 ;
    RECT 328.51 172.865 329.29 180.405 ;
    LAYER Via34 ;
    RECT 332.21 172.865 332.99 180.405 ;
    LAYER Via34 ;
    RECT 335.91 172.865 336.69 180.405 ;
    LAYER Via34 ;
    RECT 341.31 172.865 342.09 180.405 ;
    LAYER Via34 ;
    RECT 343.27 172.865 344.05 180.405 ;
    LAYER Via34 ;
    RECT 348.67 172.865 349.45 180.405 ;
    LAYER Via34 ;
    RECT 350.63 172.865 351.41 180.405 ;
    LAYER Via34 ;
    RECT 356.03 172.865 356.81 180.405 ;
    LAYER Via34 ;
    RECT 357.99 172.865 358.77 180.405 ;
    LAYER Via34 ;
    RECT 363.39 172.865 364.17 180.405 ;
    LAYER Via34 ;
    RECT 365.35 172.865 366.13 180.405 ;
    LAYER Via34 ;
    RECT 370.75 172.865 371.53 180.405 ;
    LAYER Via34 ;
    RECT 372.71 172.865 373.49 180.405 ;
    LAYER Via34 ;
    RECT 378.11 172.865 378.89 180.405 ;
    LAYER Via34 ;
    RECT 380.07 172.865 380.85 180.405 ;
    LAYER Via34 ;
    RECT 385.47 172.865 386.25 180.405 ;
    LAYER Via34 ;
    RECT 387.43 172.865 388.21 180.405 ;
    LAYER Via34 ;
    RECT 392.83 172.865 393.61 180.405 ;
    LAYER Via34 ;
    RECT 394.71 172.865 395.49 180.405 ;
    LAYER Via34 ;
    RECT 396.59 172.865 397.37 180.405 ;
    LAYER Via34 ;
    RECT 401.99 172.865 402.77 180.405 ;
    LAYER Via34 ;
    RECT 403.95 172.865 404.73 180.405 ;
    LAYER Via34 ;
    RECT 409.35 172.865 410.13 180.405 ;
    LAYER Via34 ;
    RECT 411.31 172.865 412.09 180.405 ;
    LAYER Via34 ;
    RECT 416.71 172.865 417.49 180.405 ;
    LAYER Via34 ;
    RECT 418.67 172.865 419.45 180.405 ;
    LAYER Via34 ;
    RECT 424.07 172.865 424.85 180.405 ;
    LAYER Via34 ;
    RECT 426.03 172.865 426.81 180.405 ;
    LAYER Via34 ;
    RECT 431.43 172.865 432.21 180.405 ;
    LAYER Via34 ;
    RECT 433.39 172.865 434.17 180.405 ;
    LAYER Via34 ;
    RECT 438.79 172.865 439.57 180.405 ;
    LAYER Via34 ;
    RECT 440.75 172.865 441.53 180.405 ;
    LAYER Via34 ;
    RECT 446.15 172.865 446.93 180.405 ;
    LAYER Via34 ;
    RECT 448.11 172.865 448.89 180.405 ;
    LAYER Via34 ;
    RECT 453.51 172.865 454.29 180.405 ;
    LAYER Via34 ;
    RECT 455.39 172.865 456.17 180.405 ;
    LAYER Via34 ;
    RECT 457.27 172.865 458.05 180.405 ;
    LAYER Via34 ;
    RECT 462.67 172.865 463.45 180.405 ;
    LAYER Via34 ;
    RECT 464.63 172.865 465.41 180.405 ;
    LAYER Via34 ;
    RECT 470.03 172.865 470.81 180.405 ;
    LAYER Via34 ;
    RECT 471.99 172.865 472.77 180.405 ;
    LAYER Via34 ;
    RECT 477.39 172.865 478.17 180.405 ;
    LAYER Via34 ;
    RECT 479.35 172.865 480.13 180.405 ;
    LAYER Via34 ;
    RECT 484.75 172.865 485.53 180.405 ;
    LAYER Via34 ;
    RECT 486.71 172.865 487.49 180.405 ;
    LAYER Via34 ;
    RECT 492.11 172.865 492.89 180.405 ;
    LAYER Via34 ;
    RECT 494.07 172.865 494.85 180.405 ;
    LAYER Via34 ;
    RECT 499.47 172.865 500.25 180.405 ;
    LAYER Via34 ;
    RECT 501.43 172.865 502.21 180.405 ;
    LAYER Via34 ;
    RECT 506.83 172.865 507.61 180.405 ;
    LAYER Via34 ;
    RECT 508.79 172.865 509.57 180.405 ;
    LAYER Via34 ;
    RECT 514.19 172.865 514.97 180.405 ;
    LAYER Via34 ;
    RECT 516.07 172.865 516.85 180.405 ;
    LAYER Via34 ;
    RECT 517.95 172.865 518.73 180.405 ;
    LAYER Via34 ;
    RECT 523.35 172.865 524.13 180.405 ;
    LAYER Via34 ;
    RECT 525.31 172.865 526.09 180.405 ;
    LAYER Via34 ;
    RECT 530.71 172.865 531.49 180.405 ;
    LAYER Via34 ;
    RECT 532.67 172.865 533.45 180.405 ;
    LAYER Via34 ;
    RECT 538.07 172.865 538.85 180.405 ;
    LAYER Via34 ;
    RECT 540.03 172.865 540.81 180.405 ;
    LAYER Via34 ;
    RECT 545.43 172.865 546.21 180.405 ;
    LAYER Via34 ;
    RECT 547.39 172.865 548.17 180.405 ;
    LAYER Via34 ;
    RECT 552.79 172.865 553.57 180.405 ;
    LAYER Via34 ;
    RECT 554.75 172.865 555.53 180.405 ;
    LAYER Via34 ;
    RECT 560.15 172.865 560.93 180.405 ;
    LAYER Via34 ;
    RECT 562.11 172.865 562.89 180.405 ;
    LAYER Via34 ;
    RECT 567.51 172.865 568.29 180.405 ;
    LAYER Via34 ;
    RECT 569.47 172.865 570.25 180.405 ;
    LAYER Via34 ;
    RECT 574.87 172.865 575.65 180.405 ;
    LAYER Via34 ;
    RECT 576.77 172.865 577.55 180.405 ;
    LAYER Via34 ;
    RECT 19.79 8.83 20.57 16.37 ;
    LAYER Via34 ;
    RECT 21.59 8.83 22.37 16.37 ;
    LAYER Via34 ;
    RECT 27.91 8.83 30.77 16.37 ;
    LAYER Via34 ;
    RECT 36.31 8.83 37.09 16.37 ;
    LAYER Via34 ;
    RECT 43.32 8.83 44.1 16.37 ;
    LAYER Via34 ;
    RECT 51.03 8.83 51.81 16.37 ;
    LAYER Via34 ;
    RECT 58.74 8.83 59.52 16.37 ;
    LAYER Via34 ;
    RECT 65.75 8.83 66.53 16.37 ;
    LAYER Via34 ;
    RECT 72.07 8.83 74.93 16.37 ;
    LAYER Via34 ;
    RECT 80.47 8.83 81.25 16.37 ;
    LAYER Via34 ;
    RECT 82.27 8.83 83.05 16.37 ;
    LAYER Via34 ;
    RECT 88.59 8.83 91.45 16.37 ;
    LAYER Via34 ;
    RECT 96.99 8.83 97.77 16.37 ;
    LAYER Via34 ;
    RECT 104 8.83 104.78 16.37 ;
    LAYER Via34 ;
    RECT 111.71 8.83 112.49 16.37 ;
    LAYER Via34 ;
    RECT 119.42 8.83 120.2 16.37 ;
    LAYER Via34 ;
    RECT 126.43 8.83 127.21 16.37 ;
    LAYER Via34 ;
    RECT 132.75 8.83 135.61 16.37 ;
    LAYER Via34 ;
    RECT 141.15 8.83 141.93 16.37 ;
    LAYER Via34 ;
    RECT 142.95 8.83 143.73 16.37 ;
    LAYER Via34 ;
    RECT 149.27 8.83 152.13 16.37 ;
    LAYER Via34 ;
    RECT 157.67 8.83 158.45 16.37 ;
    LAYER Via34 ;
    RECT 164.68 8.83 165.46 16.37 ;
    LAYER Via34 ;
    RECT 172.39 8.83 173.17 16.37 ;
    LAYER Via34 ;
    RECT 180.1 8.83 180.88 16.37 ;
    LAYER Via34 ;
    RECT 187.11 8.83 187.89 16.37 ;
    LAYER Via34 ;
    RECT 193.43 8.83 196.29 16.37 ;
    LAYER Via34 ;
    RECT 201.83 8.83 202.61 16.37 ;
    LAYER Via34 ;
    RECT 203.63 8.83 204.41 16.37 ;
    LAYER Via34 ;
    RECT 209.95 8.83 212.81 16.37 ;
    LAYER Via34 ;
    RECT 218.35 8.83 219.13 16.37 ;
    LAYER Via34 ;
    RECT 225.36 8.83 226.14 16.37 ;
    LAYER Via34 ;
    RECT 233.07 8.83 233.85 16.37 ;
    LAYER Via34 ;
    RECT 240.78 8.83 241.56 16.37 ;
    LAYER Via34 ;
    RECT 247.79 8.83 248.57 16.37 ;
    LAYER Via34 ;
    RECT 254.11 8.83 256.97 16.37 ;
    LAYER Via34 ;
    RECT 262.51 8.83 263.29 16.37 ;
    LAYER Via34 ;
    RECT 264.31 8.83 265.09 16.37 ;
    LAYER Via34 ;
    RECT 266.06 8.83 267.36 16.37 ;
    LAYER Via34 ;
    RECT 272.85 8.83 274.15 16.37 ;
    LAYER Via34 ;
    RECT 281.65 8.83 282.95 16.37 ;
    LAYER Via34 ;
    RECT 290.45 8.83 291.75 16.37 ;
    LAYER Via34 ;
    RECT 299.25 8.83 300.55 16.37 ;
    LAYER Via34 ;
    RECT 308.05 8.83 309.35 16.37 ;
    LAYER Via34 ;
    RECT 317.66 8.83 317.92 16.37 ;
    LAYER Via34 ;
    RECT 323.42 8.83 323.68 16.37 ;
    LAYER Via34 ;
    RECT 329.18 8.83 329.44 16.37 ;
    LAYER Via34 ;
    RECT 331.87 8.83 332.65 16.37 ;
    LAYER Via34 ;
    RECT 334.93 8.83 335.71 16.37 ;
    LAYER Via34 ;
    RECT 341.25 8.83 344.11 16.37 ;
    LAYER Via34 ;
    RECT 349.65 8.83 350.43 16.37 ;
    LAYER Via34 ;
    RECT 356.66 8.83 357.44 16.37 ;
    LAYER Via34 ;
    RECT 364.37 8.83 365.15 16.37 ;
    LAYER Via34 ;
    RECT 372.08 8.83 372.86 16.37 ;
    LAYER Via34 ;
    RECT 379.09 8.83 379.87 16.37 ;
    LAYER Via34 ;
    RECT 385.41 8.83 388.27 16.37 ;
    LAYER Via34 ;
    RECT 393.81 8.83 394.59 16.37 ;
    LAYER Via34 ;
    RECT 395.61 8.83 396.39 16.37 ;
    LAYER Via34 ;
    RECT 401.93 8.83 404.79 16.37 ;
    LAYER Via34 ;
    RECT 410.33 8.83 411.11 16.37 ;
    LAYER Via34 ;
    RECT 417.34 8.83 418.12 16.37 ;
    LAYER Via34 ;
    RECT 425.05 8.83 425.83 16.37 ;
    LAYER Via34 ;
    RECT 432.76 8.83 433.54 16.37 ;
    LAYER Via34 ;
    RECT 439.77 8.83 440.55 16.37 ;
    LAYER Via34 ;
    RECT 446.09 8.83 448.95 16.37 ;
    LAYER Via34 ;
    RECT 454.49 8.83 455.27 16.37 ;
    LAYER Via34 ;
    RECT 456.29 8.83 457.07 16.37 ;
    LAYER Via34 ;
    RECT 462.61 8.83 465.47 16.37 ;
    LAYER Via34 ;
    RECT 471.01 8.83 471.79 16.37 ;
    LAYER Via34 ;
    RECT 478.02 8.83 478.8 16.37 ;
    LAYER Via34 ;
    RECT 485.73 8.83 486.51 16.37 ;
    LAYER Via34 ;
    RECT 493.44 8.83 494.22 16.37 ;
    LAYER Via34 ;
    RECT 500.45 8.83 501.23 16.37 ;
    LAYER Via34 ;
    RECT 506.77 8.83 509.63 16.37 ;
    LAYER Via34 ;
    RECT 515.17 8.83 515.95 16.37 ;
    LAYER Via34 ;
    RECT 516.97 8.83 517.75 16.37 ;
    LAYER Via34 ;
    RECT 523.29 8.83 526.15 16.37 ;
    LAYER Via34 ;
    RECT 531.69 8.83 532.47 16.37 ;
    LAYER Via34 ;
    RECT 538.7 8.83 539.48 16.37 ;
    LAYER Via34 ;
    RECT 546.41 8.83 547.19 16.37 ;
    LAYER Via34 ;
    RECT 554.12 8.83 554.9 16.37 ;
    LAYER Via34 ;
    RECT 561.13 8.83 561.91 16.37 ;
    LAYER Via34 ;
    RECT 567.45 8.83 570.31 16.37 ;
    LAYER Via34 ;
    RECT 575.85 8.83 576.63 16.37 ;
    LAYER Via34 ;
    RECT 577.65 8.83 578.43 16.37 ;
    LAYER Via34 ;
    RECT 581.85 29.025 589.39 29.805 ;
    LAYER Via34 ;
    RECT 581.85 54.855 589.39 57.195 ;
    LAYER Via34 ;
    RECT 581.85 63.36 589.39 67.78 ;
    LAYER Via34 ;
    RECT 581.85 74.435 589.39 74.695 ;
    LAYER Via34 ;
    RECT 581.85 87.195 589.39 89.015 ;
    LAYER Via34 ;
    RECT 581.85 121.125 589.39 121.905 ;
    LAYER Via34 ;
    RECT 581.85 126.185 589.39 126.965 ;
    LAYER Via34 ;
    RECT 581.85 131.245 589.39 132.025 ;
    LAYER Via34 ;
    RECT 581.85 136.305 589.39 137.085 ;
    LAYER Via34 ;
    RECT 581.85 141.365 589.39 142.145 ;
    LAYER Via34 ;
    RECT 581.85 146.425 589.39 147.205 ;
    LAYER Via34 ;
    RECT 581.85 151.485 589.39 152.265 ;
    LAYER Via34 ;
    RECT 581.85 156.545 589.39 157.325 ;
    LAYER Via34 ;
    RECT 581.85 161.605 589.39 162.385 ;
    LAYER Via34 ;
    RECT 581.85 166.665 589.39 167.445 ;
    LAYER Via34 ;
    RECT 581.85 170.115 589.39 170.895 ;
    LAYER Via34 ;
    RECT 8.83 29.025 16.37 29.805 ;
    LAYER Via34 ;
    RECT 8.83 54.855 16.37 57.195 ;
    LAYER Via34 ;
    RECT 8.83 63.36 16.37 67.78 ;
    LAYER Via34 ;
    RECT 8.83 74.435 16.37 74.695 ;
    LAYER Via34 ;
    RECT 8.83 87.195 16.37 89.015 ;
    LAYER Via34 ;
    RECT 8.83 121.125 16.37 121.905 ;
    LAYER Via34 ;
    RECT 8.83 126.185 16.37 126.965 ;
    LAYER Via34 ;
    RECT 8.83 131.245 16.37 132.025 ;
    LAYER Via34 ;
    RECT 8.83 136.305 16.37 137.085 ;
    LAYER Via34 ;
    RECT 8.83 141.365 16.37 142.145 ;
    LAYER Via34 ;
    RECT 8.83 146.425 16.37 147.205 ;
    LAYER Via34 ;
    RECT 8.83 151.485 16.37 152.265 ;
    LAYER Via34 ;
    RECT 8.83 156.545 16.37 157.325 ;
    LAYER Via34 ;
    RECT 8.83 161.605 16.37 162.385 ;
    LAYER Via34 ;
    RECT 8.83 166.665 16.37 167.445 ;
    LAYER Via34 ;
    RECT 8.83 170.115 16.37 170.895 ;
    END
  #BEGINEXT "VSI SIGNATURE 1.0"
    #CREATOR "Artisan Components, Inc." ;
    #DATE "2001-04-10" ;
    #REVISION "1.0" ;
    #ENDEXT
  END ram_256x16A

MACRO rom_512x16A
  CLASS RING ;
  FOREIGN rom_512x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 368.165 BY 186.845 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 88.705 21.2 89.805 22.3 ;
      LAYER Metal2 ;
      RECT 88.705 21.2 89.805 22.3 ;
      LAYER Metal3 ;
      RECT 88.705 21.2 89.805 22.3 ;
      LAYER Metal4 ;
      RECT 88.705 21.2 89.805 22.3 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 84.205 21.2 85.305 22.3 ;
      LAYER Metal2 ;
      RECT 84.205 21.2 85.305 22.3 ;
      LAYER Metal3 ;
      RECT 84.205 21.2 85.305 22.3 ;
      LAYER Metal4 ;
      RECT 84.205 21.2 85.305 22.3 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 79.705 21.2 80.805 22.3 ;
      LAYER Metal2 ;
      RECT 79.705 21.2 80.805 22.3 ;
      LAYER Metal3 ;
      RECT 79.705 21.2 80.805 22.3 ;
      LAYER Metal4 ;
      RECT 79.705 21.2 80.805 22.3 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 70.705 21.2 71.805 22.3 ;
      LAYER Metal2 ;
      RECT 70.705 21.2 71.805 22.3 ;
      LAYER Metal3 ;
      RECT 70.705 21.2 71.805 22.3 ;
      LAYER Metal4 ;
      RECT 70.705 21.2 71.805 22.3 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 61.705 21.2 62.805 22.3 ;
      LAYER Metal2 ;
      RECT 61.705 21.2 62.805 22.3 ;
      LAYER Metal3 ;
      RECT 61.705 21.2 62.805 22.3 ;
      LAYER Metal4 ;
      RECT 61.705 21.2 62.805 22.3 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 57.205 21.2 58.305 22.3 ;
      LAYER Metal2 ;
      RECT 57.205 21.2 58.305 22.3 ;
      LAYER Metal3 ;
      RECT 57.205 21.2 58.305 22.3 ;
      LAYER Metal4 ;
      RECT 57.205 21.2 58.305 22.3 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 52.705 21.2 53.805 22.3 ;
      LAYER Metal2 ;
      RECT 52.705 21.2 53.805 22.3 ;
      LAYER Metal3 ;
      RECT 52.705 21.2 53.805 22.3 ;
      LAYER Metal4 ;
      RECT 52.705 21.2 53.805 22.3 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 43.705 21.2 44.805 22.3 ;
      LAYER Metal2 ;
      RECT 43.705 21.2 44.805 22.3 ;
      LAYER Metal3 ;
      RECT 43.705 21.2 44.805 22.3 ;
      LAYER Metal4 ;
      RECT 43.705 21.2 44.805 22.3 ;
      END
    END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 39.205 21.2 40.305 22.3 ;
      LAYER Metal2 ;
      RECT 39.205 21.2 40.305 22.3 ;
      LAYER Metal3 ;
      RECT 39.205 21.2 40.305 22.3 ;
      LAYER Metal4 ;
      RECT 39.205 21.2 40.305 22.3 ;
      END
    END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 112.02 21.2 113.12 22.3 ;
      LAYER Metal2 ;
      RECT 112.02 21.2 113.12 22.3 ;
      LAYER Metal3 ;
      RECT 112.02 21.2 113.12 22.3 ;
      LAYER Metal4 ;
      RECT 112.02 21.2 113.12 22.3 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    AntennaGateArea  0.792 ;
    PORT
      LAYER Metal1 ;
      RECT 110.32 21.2 111.42 22.3 ;
      LAYER Metal2 ;
      RECT 110.32 21.2 111.42 22.3 ;
      LAYER Metal3 ;
      RECT 110.32 21.2 111.42 22.3 ;
      LAYER Metal4 ;
      RECT 110.32 21.2 111.42 22.3 ;
      END
    END CLK
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 141.575 21.2 142.675 22.3 ;
      LAYER Metal2 ;
      RECT 141.575 21.2 142.675 22.3 ;
      LAYER Metal3 ;
      RECT 141.575 21.2 142.675 22.3 ;
      LAYER Metal4 ;
      RECT 141.575 21.2 142.675 22.3 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 275.475 21.2 276.575 22.3 ;
      LAYER Metal2 ;
      RECT 275.475 21.2 276.575 22.3 ;
      LAYER Metal3 ;
      RECT 275.475 21.2 276.575 22.3 ;
      LAYER Metal4 ;
      RECT 275.475 21.2 276.575 22.3 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 278.535 21.2 279.635 22.3 ;
      LAYER Metal2 ;
      RECT 278.535 21.2 279.635 22.3 ;
      LAYER Metal3 ;
      RECT 278.535 21.2 279.635 22.3 ;
      LAYER Metal4 ;
      RECT 278.535 21.2 279.635 22.3 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 302.255 21.2 303.355 22.3 ;
      LAYER Metal2 ;
      RECT 302.255 21.2 303.355 22.3 ;
      LAYER Metal3 ;
      RECT 302.255 21.2 303.355 22.3 ;
      LAYER Metal4 ;
      RECT 302.255 21.2 303.355 22.3 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 305.315 21.2 306.415 22.3 ;
      LAYER Metal2 ;
      RECT 305.315 21.2 306.415 22.3 ;
      LAYER Metal3 ;
      RECT 305.315 21.2 306.415 22.3 ;
      LAYER Metal4 ;
      RECT 305.315 21.2 306.415 22.3 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 329.035 21.2 330.135 22.3 ;
      LAYER Metal2 ;
      RECT 329.035 21.2 330.135 22.3 ;
      LAYER Metal3 ;
      RECT 329.035 21.2 330.135 22.3 ;
      LAYER Metal4 ;
      RECT 329.035 21.2 330.135 22.3 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 332.095 21.2 333.195 22.3 ;
      LAYER Metal2 ;
      RECT 332.095 21.2 333.195 22.3 ;
      LAYER Metal3 ;
      RECT 332.095 21.2 333.195 22.3 ;
      LAYER Metal4 ;
      RECT 332.095 21.2 333.195 22.3 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 144.635 21.2 145.735 22.3 ;
      LAYER Metal2 ;
      RECT 144.635 21.2 145.735 22.3 ;
      LAYER Metal3 ;
      RECT 144.635 21.2 145.735 22.3 ;
      LAYER Metal4 ;
      RECT 144.635 21.2 145.735 22.3 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 168.355 21.2 169.455 22.3 ;
      LAYER Metal2 ;
      RECT 168.355 21.2 169.455 22.3 ;
      LAYER Metal3 ;
      RECT 168.355 21.2 169.455 22.3 ;
      LAYER Metal4 ;
      RECT 168.355 21.2 169.455 22.3 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 171.415 21.2 172.515 22.3 ;
      LAYER Metal2 ;
      RECT 171.415 21.2 172.515 22.3 ;
      LAYER Metal3 ;
      RECT 171.415 21.2 172.515 22.3 ;
      LAYER Metal4 ;
      RECT 171.415 21.2 172.515 22.3 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 195.135 21.2 196.235 22.3 ;
      LAYER Metal2 ;
      RECT 195.135 21.2 196.235 22.3 ;
      LAYER Metal3 ;
      RECT 195.135 21.2 196.235 22.3 ;
      LAYER Metal4 ;
      RECT 195.135 21.2 196.235 22.3 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 198.195 21.2 199.295 22.3 ;
      LAYER Metal2 ;
      RECT 198.195 21.2 199.295 22.3 ;
      LAYER Metal3 ;
      RECT 198.195 21.2 199.295 22.3 ;
      LAYER Metal4 ;
      RECT 198.195 21.2 199.295 22.3 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 221.915 21.2 223.015 22.3 ;
      LAYER Metal2 ;
      RECT 221.915 21.2 223.015 22.3 ;
      LAYER Metal3 ;
      RECT 221.915 21.2 223.015 22.3 ;
      LAYER Metal4 ;
      RECT 221.915 21.2 223.015 22.3 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 224.975 21.2 226.075 22.3 ;
      LAYER Metal2 ;
      RECT 224.975 21.2 226.075 22.3 ;
      LAYER Metal3 ;
      RECT 224.975 21.2 226.075 22.3 ;
      LAYER Metal4 ;
      RECT 224.975 21.2 226.075 22.3 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 248.695 21.2 249.795 22.3 ;
      LAYER Metal2 ;
      RECT 248.695 21.2 249.795 22.3 ;
      LAYER Metal3 ;
      RECT 248.695 21.2 249.795 22.3 ;
      LAYER Metal4 ;
      RECT 248.695 21.2 249.795 22.3 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 251.755 21.2 252.855 22.3 ;
      LAYER Metal2 ;
      RECT 251.755 21.2 252.855 22.3 ;
      LAYER Metal3 ;
      RECT 251.755 21.2 252.855 22.3 ;
      LAYER Metal4 ;
      RECT 251.755 21.2 252.855 22.3 ;
      END
    END Q[9]
  PIN VDD
    DIRECTION OUTPUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 368.165 176.845 0 186.845 ;
      LAYER Metal5 ;
      RECT 0 0 368.165 10 ;
      LAYER Metal3 ;
      RECT 368.165 176.845 0 186.845 ;
      LAYER Metal3 ;
      RECT 0 0 368.165 10 ;
      LAYER Metal4 ;
      RECT 358.165 0 368.165 186.845 ;
      LAYER Metal4 ;
      RECT 0 186.845 10 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION OUTPUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 357.565 166.245 10.6 176.245 ;
      LAYER Metal5 ;
      RECT 10.6 10.6 357.565 20.6 ;
      LAYER Metal3 ;
      RECT 357.565 166.245 10.6 176.245 ;
      LAYER Metal3 ;
      RECT 10.6 10.6 357.565 20.6 ;
      LAYER Metal4 ;
      RECT 347.565 10.6 357.565 176.245 ;
      LAYER Metal4 ;
      RECT 10.6 176.245 20.6 10.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Metal1 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Metal2 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Metal3 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Metal4 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Via12 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Via23 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Via34 ;
    RECT 21.2 21.2 346.965 165.645 ;
    LAYER Via34 ;
    RECT 347.755 166.435 357.375 176.055 ;
    LAYER Via34 ;
    RECT 10.79 10.79 20.41 20.41 ;
    LAYER Via34 ;
    RECT 347.755 10.79 357.375 20.41 ;
    LAYER Via34 ;
    RECT 10.79 166.435 20.41 176.055 ;
    LAYER Via34 ;
    RECT 358.355 177.035 367.975 186.655 ;
    LAYER Via34 ;
    RECT 0.19 0.19 9.81 9.81 ;
    LAYER Via34 ;
    RECT 358.355 0.19 367.975 9.81 ;
    LAYER Via34 ;
    RECT 0.19 177.035 9.81 186.655 ;
    LAYER Metal4 ;
    RECT 25.445 165.645 26.445 186.845 ;
    LAYER Metal4 ;
    RECT 29.105 165.645 37.605 186.845 ;
    LAYER Metal4 ;
    RECT 47.805 165.645 56.805 186.845 ;
    LAYER Metal4 ;
    RECT 67.005 165.645 76.005 186.845 ;
    LAYER Metal4 ;
    RECT 86.205 165.645 95.205 186.845 ;
    LAYER Metal4 ;
    RECT 99.32 165.645 101.92 186.845 ;
    LAYER Metal4 ;
    RECT 106.76 165.645 110.56 186.845 ;
    LAYER Metal4 ;
    RECT 115.4 165.645 119.2 186.845 ;
    LAYER Metal4 ;
    RECT 124.01 165.645 127.31 186.845 ;
    LAYER Metal4 ;
    RECT 27.505 21.2 29.505 0 ;
    LAYER Metal4 ;
    RECT 36.505 21.2 38.505 0 ;
    LAYER Metal4 ;
    RECT 45.505 21.2 47.505 0 ;
    LAYER Metal4 ;
    RECT 54.505 21.2 56.505 0 ;
    LAYER Metal4 ;
    RECT 63.505 21.2 65.505 0 ;
    LAYER Metal4 ;
    RECT 72.505 21.2 74.505 0 ;
    LAYER Metal4 ;
    RECT 81.505 21.2 83.505 0 ;
    LAYER Metal4 ;
    RECT 90.505 21.2 92.505 0 ;
    LAYER Metal4 ;
    RECT 100.02 21.2 108.02 0 ;
    LAYER Metal4 ;
    RECT 124.01 21.2 127.31 0 ;
    LAYER Metal4 ;
    RECT 129.765 21.2 130.765 0 ;
    LAYER Metal4 ;
    RECT 132.685 21.2 133.685 0 ;
    LAYER Metal4 ;
    RECT 135.605 21.2 136.605 0 ;
    LAYER Metal4 ;
    RECT 138.525 21.2 139.525 0 ;
    LAYER Metal4 ;
    RECT 147.785 21.2 148.785 0 ;
    LAYER Metal4 ;
    RECT 150.705 21.2 151.705 0 ;
    LAYER Metal4 ;
    RECT 153.625 21.2 154.625 0 ;
    LAYER Metal4 ;
    RECT 156.545 21.2 157.545 0 ;
    LAYER Metal4 ;
    RECT 159.465 21.2 160.465 0 ;
    LAYER Metal4 ;
    RECT 162.385 21.2 163.385 0 ;
    LAYER Metal4 ;
    RECT 165.305 21.2 166.305 0 ;
    LAYER Metal4 ;
    RECT 174.565 21.2 175.565 0 ;
    LAYER Metal4 ;
    RECT 177.485 21.2 178.485 0 ;
    LAYER Metal4 ;
    RECT 180.405 21.2 181.405 0 ;
    LAYER Metal4 ;
    RECT 183.325 21.2 184.325 0 ;
    LAYER Metal4 ;
    RECT 186.245 21.2 187.245 0 ;
    LAYER Metal4 ;
    RECT 189.165 21.2 190.165 0 ;
    LAYER Metal4 ;
    RECT 192.085 21.2 193.085 0 ;
    LAYER Metal4 ;
    RECT 201.345 21.2 202.345 0 ;
    LAYER Metal4 ;
    RECT 204.265 21.2 205.265 0 ;
    LAYER Metal4 ;
    RECT 207.185 21.2 208.185 0 ;
    LAYER Metal4 ;
    RECT 210.105 21.2 211.105 0 ;
    LAYER Metal4 ;
    RECT 213.025 21.2 214.025 0 ;
    LAYER Metal4 ;
    RECT 215.945 21.2 216.945 0 ;
    LAYER Metal4 ;
    RECT 218.865 21.2 219.865 0 ;
    LAYER Metal4 ;
    RECT 228.125 21.2 229.125 0 ;
    LAYER Metal4 ;
    RECT 231.045 21.2 232.045 0 ;
    LAYER Metal4 ;
    RECT 233.965 21.2 234.965 0 ;
    LAYER Metal4 ;
    RECT 236.885 21.2 237.885 0 ;
    LAYER Metal4 ;
    RECT 239.805 21.2 240.805 0 ;
    LAYER Metal4 ;
    RECT 242.725 21.2 243.725 0 ;
    LAYER Metal4 ;
    RECT 245.645 21.2 246.645 0 ;
    LAYER Metal4 ;
    RECT 254.905 21.2 255.905 0 ;
    LAYER Metal4 ;
    RECT 257.825 21.2 258.825 0 ;
    LAYER Metal4 ;
    RECT 260.745 21.2 261.745 0 ;
    LAYER Metal4 ;
    RECT 263.665 21.2 264.665 0 ;
    LAYER Metal4 ;
    RECT 266.585 21.2 267.585 0 ;
    LAYER Metal4 ;
    RECT 269.505 21.2 270.505 0 ;
    LAYER Metal4 ;
    RECT 272.425 21.2 273.425 0 ;
    LAYER Metal4 ;
    RECT 281.685 21.2 282.685 0 ;
    LAYER Metal4 ;
    RECT 284.605 21.2 285.605 0 ;
    LAYER Metal4 ;
    RECT 287.525 21.2 288.525 0 ;
    LAYER Metal4 ;
    RECT 290.445 21.2 291.445 0 ;
    LAYER Metal4 ;
    RECT 293.365 21.2 294.365 0 ;
    LAYER Metal4 ;
    RECT 296.285 21.2 297.285 0 ;
    LAYER Metal4 ;
    RECT 299.205 21.2 300.205 0 ;
    LAYER Metal4 ;
    RECT 308.465 21.2 309.465 0 ;
    LAYER Metal4 ;
    RECT 311.385 21.2 312.385 0 ;
    LAYER Metal4 ;
    RECT 314.305 21.2 315.305 0 ;
    LAYER Metal4 ;
    RECT 317.225 21.2 318.225 0 ;
    LAYER Metal4 ;
    RECT 320.145 21.2 321.145 0 ;
    LAYER Metal4 ;
    RECT 323.065 21.2 324.065 0 ;
    LAYER Metal4 ;
    RECT 325.985 21.2 326.985 0 ;
    LAYER Metal4 ;
    RECT 335.245 21.2 336.245 0 ;
    LAYER Metal4 ;
    RECT 338.165 21.2 339.165 0 ;
    LAYER Metal4 ;
    RECT 341.085 21.2 342.085 0 ;
    LAYER Metal4 ;
    RECT 344.005 21.2 345.005 0 ;
    LAYER Metal3 ;
    RECT 346.965 23.7 368.165 24.7 ;
    LAYER Metal3 ;
    RECT 346.965 47.04 368.165 49.04 ;
    LAYER Metal3 ;
    RECT 346.965 54.64 368.165 56.14 ;
    LAYER Metal3 ;
    RECT 346.965 58.7 368.165 60.7 ;
    LAYER Metal3 ;
    RECT 346.965 70.5 368.165 72.5 ;
    LAYER Metal3 ;
    RECT 346.965 78.41 368.165 79.31 ;
    LAYER Metal3 ;
    RECT 346.965 86.38 368.165 87.78 ;
    LAYER Metal3 ;
    RECT 346.965 90.375 368.165 91.575 ;
    LAYER Metal3 ;
    RECT 346.965 97.63 368.165 99.63 ;
    LAYER Metal3 ;
    RECT 346.965 109.235 368.165 111.235 ;
    LAYER Metal3 ;
    RECT 346.965 113.755 368.165 115.255 ;
    LAYER Metal3 ;
    RECT 346.965 120.715 368.165 122.715 ;
    LAYER Metal3 ;
    RECT 346.965 125.085 368.165 127.885 ;
    LAYER Metal3 ;
    RECT 21.2 24.675 0 25.675 ;
    LAYER Metal3 ;
    RECT 21.2 39.14 0 44.14 ;
    LAYER Metal3 ;
    RECT 21.2 56.5 0 63.5 ;
    LAYER Metal3 ;
    RECT 21.2 77.86 0 78.86 ;
    LAYER Metal3 ;
    RECT 21.2 88.25 0 89.85 ;
    LAYER Metal3 ;
    RECT 21.2 97.63 0 99.63 ;
    LAYER Metal3 ;
    RECT 21.2 109.81 0 112.81 ;
    LAYER Metal3 ;
    RECT 21.2 120.215 0 123.215 ;
    LAYER Metal4 ;
    RECT 23.305 165.645 24.785 176.245 ;
    LAYER Metal4 ;
    RECT 27.225 165.645 28.225 176.245 ;
    LAYER Metal4 ;
    RECT 38.205 165.645 47.205 176.245 ;
    LAYER Metal4 ;
    RECT 57.405 165.645 66.405 176.245 ;
    LAYER Metal4 ;
    RECT 76.605 165.645 85.605 176.245 ;
    LAYER Metal4 ;
    RECT 95.86 165.645 98.86 176.245 ;
    LAYER Metal4 ;
    RECT 102.44 165.645 106.24 176.245 ;
    LAYER Metal4 ;
    RECT 111.08 165.645 114.88 176.245 ;
    LAYER Metal4 ;
    RECT 119.72 165.645 122.32 176.245 ;
    LAYER Metal4 ;
    RECT 127.795 165.645 129.295 176.245 ;
    LAYER Metal4 ;
    RECT 131.185 165.645 135.185 176.245 ;
    LAYER Metal4 ;
    RECT 137.025 165.645 141.025 176.245 ;
    LAYER Metal4 ;
    RECT 142.455 165.645 144.855 176.245 ;
    LAYER Metal4 ;
    RECT 146.285 165.645 150.285 176.245 ;
    LAYER Metal4 ;
    RECT 152.125 165.645 156.125 176.245 ;
    LAYER Metal4 ;
    RECT 157.965 165.645 161.965 176.245 ;
    LAYER Metal4 ;
    RECT 163.805 165.645 167.805 176.245 ;
    LAYER Metal4 ;
    RECT 169.235 165.645 171.635 176.245 ;
    LAYER Metal4 ;
    RECT 173.065 165.645 177.065 176.245 ;
    LAYER Metal4 ;
    RECT 178.905 165.645 182.905 176.245 ;
    LAYER Metal4 ;
    RECT 184.745 165.645 188.745 176.245 ;
    LAYER Metal4 ;
    RECT 190.585 165.645 194.585 176.245 ;
    LAYER Metal4 ;
    RECT 196.015 165.645 198.415 176.245 ;
    LAYER Metal4 ;
    RECT 199.845 165.645 203.845 176.245 ;
    LAYER Metal4 ;
    RECT 205.685 165.645 209.685 176.245 ;
    LAYER Metal4 ;
    RECT 211.525 165.645 215.525 176.245 ;
    LAYER Metal4 ;
    RECT 217.365 165.645 221.365 176.245 ;
    LAYER Metal4 ;
    RECT 222.795 165.645 225.195 176.245 ;
    LAYER Metal4 ;
    RECT 226.625 165.645 230.625 176.245 ;
    LAYER Metal4 ;
    RECT 232.465 165.645 236.465 176.245 ;
    LAYER Metal4 ;
    RECT 238.305 165.645 242.305 176.245 ;
    LAYER Metal4 ;
    RECT 244.145 165.645 248.145 176.245 ;
    LAYER Metal4 ;
    RECT 249.575 165.645 251.975 176.245 ;
    LAYER Metal4 ;
    RECT 253.405 165.645 257.405 176.245 ;
    LAYER Metal4 ;
    RECT 259.245 165.645 263.245 176.245 ;
    LAYER Metal4 ;
    RECT 265.085 165.645 269.085 176.245 ;
    LAYER Metal4 ;
    RECT 270.925 165.645 274.925 176.245 ;
    LAYER Metal4 ;
    RECT 276.355 165.645 278.755 176.245 ;
    LAYER Metal4 ;
    RECT 280.185 165.645 284.185 176.245 ;
    LAYER Metal4 ;
    RECT 286.025 165.645 290.025 176.245 ;
    LAYER Metal4 ;
    RECT 291.865 165.645 295.865 176.245 ;
    LAYER Metal4 ;
    RECT 297.705 165.645 301.705 176.245 ;
    LAYER Metal4 ;
    RECT 303.135 165.645 305.535 176.245 ;
    LAYER Metal4 ;
    RECT 306.965 165.645 310.965 176.245 ;
    LAYER Metal4 ;
    RECT 312.805 165.645 316.805 176.245 ;
    LAYER Metal4 ;
    RECT 318.645 165.645 322.645 176.245 ;
    LAYER Metal4 ;
    RECT 324.485 165.645 328.485 176.245 ;
    LAYER Metal4 ;
    RECT 329.915 165.645 332.315 176.245 ;
    LAYER Metal4 ;
    RECT 333.745 165.645 337.745 176.245 ;
    LAYER Metal4 ;
    RECT 339.585 165.645 343.585 176.245 ;
    LAYER Metal4 ;
    RECT 344.505 165.645 345.045 176.245 ;
    LAYER Metal4 ;
    RECT 23.3 21.2 24.8 10.6 ;
    LAYER Metal4 ;
    RECT 31.005 21.2 35.005 10.6 ;
    LAYER Metal4 ;
    RECT 41.005 21.2 43.005 10.6 ;
    LAYER Metal4 ;
    RECT 50.005 21.2 52.005 10.6 ;
    LAYER Metal4 ;
    RECT 59.005 21.2 61.005 10.6 ;
    LAYER Metal4 ;
    RECT 68.005 21.2 70.005 10.6 ;
    LAYER Metal4 ;
    RECT 77.005 21.2 79.005 10.6 ;
    LAYER Metal4 ;
    RECT 86.005 21.2 88.005 10.6 ;
    LAYER Metal4 ;
    RECT 95.86 21.2 98.86 10.6 ;
    LAYER Metal4 ;
    RECT 113.82 21.2 121.82 10.6 ;
    LAYER Metal4 ;
    RECT 127.795 21.2 129.295 10.6 ;
    LAYER Metal4 ;
    RECT 131.225 21.2 132.225 10.6 ;
    LAYER Metal4 ;
    RECT 134.145 21.2 135.145 10.6 ;
    LAYER Metal4 ;
    RECT 137.065 21.2 138.065 10.6 ;
    LAYER Metal4 ;
    RECT 139.985 21.2 140.985 10.6 ;
    LAYER Metal4 ;
    RECT 143.155 21.2 144.155 10.6 ;
    LAYER Metal4 ;
    RECT 146.325 21.2 147.325 10.6 ;
    LAYER Metal4 ;
    RECT 149.245 21.2 150.245 10.6 ;
    LAYER Metal4 ;
    RECT 152.165 21.2 153.165 10.6 ;
    LAYER Metal4 ;
    RECT 155.085 21.2 156.085 10.6 ;
    LAYER Metal4 ;
    RECT 158.005 21.2 159.005 10.6 ;
    LAYER Metal4 ;
    RECT 160.925 21.2 161.925 10.6 ;
    LAYER Metal4 ;
    RECT 163.845 21.2 164.845 10.6 ;
    LAYER Metal4 ;
    RECT 166.765 21.2 167.765 10.6 ;
    LAYER Metal4 ;
    RECT 169.935 21.2 170.935 10.6 ;
    LAYER Metal4 ;
    RECT 173.105 21.2 174.105 10.6 ;
    LAYER Metal4 ;
    RECT 176.025 21.2 177.025 10.6 ;
    LAYER Metal4 ;
    RECT 178.945 21.2 179.945 10.6 ;
    LAYER Metal4 ;
    RECT 181.865 21.2 182.865 10.6 ;
    LAYER Metal4 ;
    RECT 184.785 21.2 185.785 10.6 ;
    LAYER Metal4 ;
    RECT 187.705 21.2 188.705 10.6 ;
    LAYER Metal4 ;
    RECT 190.625 21.2 191.625 10.6 ;
    LAYER Metal4 ;
    RECT 193.545 21.2 194.545 10.6 ;
    LAYER Metal4 ;
    RECT 196.715 21.2 197.715 10.6 ;
    LAYER Metal4 ;
    RECT 199.885 21.2 200.885 10.6 ;
    LAYER Metal4 ;
    RECT 202.805 21.2 203.805 10.6 ;
    LAYER Metal4 ;
    RECT 205.725 21.2 206.725 10.6 ;
    LAYER Metal4 ;
    RECT 208.645 21.2 209.645 10.6 ;
    LAYER Metal4 ;
    RECT 211.565 21.2 212.565 10.6 ;
    LAYER Metal4 ;
    RECT 214.485 21.2 215.485 10.6 ;
    LAYER Metal4 ;
    RECT 217.405 21.2 218.405 10.6 ;
    LAYER Metal4 ;
    RECT 220.325 21.2 221.325 10.6 ;
    LAYER Metal4 ;
    RECT 223.495 21.2 224.495 10.6 ;
    LAYER Metal4 ;
    RECT 226.665 21.2 227.665 10.6 ;
    LAYER Metal4 ;
    RECT 229.585 21.2 230.585 10.6 ;
    LAYER Metal4 ;
    RECT 232.505 21.2 233.505 10.6 ;
    LAYER Metal4 ;
    RECT 235.425 21.2 236.425 10.6 ;
    LAYER Metal4 ;
    RECT 238.345 21.2 239.345 10.6 ;
    LAYER Metal4 ;
    RECT 241.265 21.2 242.265 10.6 ;
    LAYER Metal4 ;
    RECT 244.185 21.2 245.185 10.6 ;
    LAYER Metal4 ;
    RECT 247.105 21.2 248.105 10.6 ;
    LAYER Metal4 ;
    RECT 250.275 21.2 251.275 10.6 ;
    LAYER Metal4 ;
    RECT 253.445 21.2 254.445 10.6 ;
    LAYER Metal4 ;
    RECT 256.365 21.2 257.365 10.6 ;
    LAYER Metal4 ;
    RECT 259.285 21.2 260.285 10.6 ;
    LAYER Metal4 ;
    RECT 262.205 21.2 263.205 10.6 ;
    LAYER Metal4 ;
    RECT 265.125 21.2 266.125 10.6 ;
    LAYER Metal4 ;
    RECT 268.045 21.2 269.045 10.6 ;
    LAYER Metal4 ;
    RECT 270.965 21.2 271.965 10.6 ;
    LAYER Metal4 ;
    RECT 273.885 21.2 274.885 10.6 ;
    LAYER Metal4 ;
    RECT 277.055 21.2 278.055 10.6 ;
    LAYER Metal4 ;
    RECT 280.225 21.2 281.225 10.6 ;
    LAYER Metal4 ;
    RECT 283.145 21.2 284.145 10.6 ;
    LAYER Metal4 ;
    RECT 286.065 21.2 287.065 10.6 ;
    LAYER Metal4 ;
    RECT 288.985 21.2 289.985 10.6 ;
    LAYER Metal4 ;
    RECT 291.905 21.2 292.905 10.6 ;
    LAYER Metal4 ;
    RECT 294.825 21.2 295.825 10.6 ;
    LAYER Metal4 ;
    RECT 297.745 21.2 298.745 10.6 ;
    LAYER Metal4 ;
    RECT 300.665 21.2 301.665 10.6 ;
    LAYER Metal4 ;
    RECT 303.835 21.2 304.835 10.6 ;
    LAYER Metal4 ;
    RECT 307.005 21.2 308.005 10.6 ;
    LAYER Metal4 ;
    RECT 309.925 21.2 310.925 10.6 ;
    LAYER Metal4 ;
    RECT 312.845 21.2 313.845 10.6 ;
    LAYER Metal4 ;
    RECT 315.765 21.2 316.765 10.6 ;
    LAYER Metal4 ;
    RECT 318.685 21.2 319.685 10.6 ;
    LAYER Metal4 ;
    RECT 321.605 21.2 322.605 10.6 ;
    LAYER Metal4 ;
    RECT 324.525 21.2 325.525 10.6 ;
    LAYER Metal4 ;
    RECT 327.445 21.2 328.445 10.6 ;
    LAYER Metal4 ;
    RECT 330.615 21.2 331.615 10.6 ;
    LAYER Metal4 ;
    RECT 333.785 21.2 334.785 10.6 ;
    LAYER Metal4 ;
    RECT 336.705 21.2 337.705 10.6 ;
    LAYER Metal4 ;
    RECT 339.625 21.2 340.625 10.6 ;
    LAYER Metal4 ;
    RECT 342.545 21.2 343.545 10.6 ;
    LAYER Metal3 ;
    RECT 346.965 25.585 357.565 26.585 ;
    LAYER Metal3 ;
    RECT 346.965 42.64 357.565 44.84 ;
    LAYER Metal3 ;
    RECT 346.965 49.56 357.565 51.56 ;
    LAYER Metal3 ;
    RECT 346.965 68.115 357.565 69.535 ;
    LAYER Metal3 ;
    RECT 346.965 72.96 357.565 73.92 ;
    LAYER Metal3 ;
    RECT 346.965 79.83 357.565 80.73 ;
    LAYER Metal3 ;
    RECT 346.965 88.25 357.565 89.75 ;
    LAYER Metal3 ;
    RECT 346.965 96.21 357.565 97.17 ;
    LAYER Metal3 ;
    RECT 346.965 100.16 357.565 101.58 ;
    LAYER Metal3 ;
    RECT 346.965 116.995 357.565 119.995 ;
    LAYER Metal3 ;
    RECT 346.965 134.305 357.565 136.825 ;
    LAYER Metal3 ;
    RECT 346.965 137.565 357.565 140.085 ;
    LAYER Metal3 ;
    RECT 346.965 140.825 357.565 143.345 ;
    LAYER Metal3 ;
    RECT 346.965 144.085 357.565 146.605 ;
    LAYER Metal3 ;
    RECT 346.965 147.345 357.565 149.865 ;
    LAYER Metal3 ;
    RECT 346.965 150.605 357.565 153.125 ;
    LAYER Metal3 ;
    RECT 346.965 153.865 357.565 156.385 ;
    LAYER Metal3 ;
    RECT 346.965 157.125 357.565 159.645 ;
    LAYER Metal3 ;
    RECT 346.965 161.195 357.565 163.715 ;
    LAYER Metal3 ;
    RECT 21.2 30.59 10.6 35.59 ;
    LAYER Metal3 ;
    RECT 21.2 46.34 10.6 49.34 ;
    LAYER Metal3 ;
    RECT 21.2 64.14 10.6 67.64 ;
    LAYER Metal3 ;
    RECT 21.2 72.885 10.6 73.885 ;
    LAYER Metal3 ;
    RECT 21.2 79.78 10.6 80.78 ;
    LAYER Metal3 ;
    RECT 21.2 86.53 10.6 87.65 ;
    LAYER Metal3 ;
    RECT 21.2 95.705 10.6 97.105 ;
    LAYER Metal3 ;
    RECT 21.2 105.02 10.6 108.02 ;
    LAYER Metal3 ;
    RECT 21.2 124.655 10.6 127.655 ;
    LAYER Via34 ;
    RECT 25.555 177.035 26.335 186.655 ;
    LAYER Via34 ;
    RECT 29.325 177.035 37.385 186.655 ;
    LAYER Via34 ;
    RECT 48.015 177.035 56.595 186.655 ;
    LAYER Via34 ;
    RECT 67.215 177.035 75.795 186.655 ;
    LAYER Via34 ;
    RECT 86.415 177.035 94.995 186.655 ;
    LAYER Via34 ;
    RECT 99.45 177.035 101.79 186.655 ;
    LAYER Via34 ;
    RECT 106.97 177.035 110.35 186.655 ;
    LAYER Via34 ;
    RECT 115.61 177.035 118.99 186.655 ;
    LAYER Via34 ;
    RECT 124.23 177.035 127.09 186.655 ;
    LAYER Via34 ;
    RECT 27.595 0.19 29.415 9.81 ;
    LAYER Via34 ;
    RECT 36.595 0.19 38.415 9.81 ;
    LAYER Via34 ;
    RECT 45.595 0.19 47.415 9.81 ;
    LAYER Via34 ;
    RECT 54.595 0.19 56.415 9.81 ;
    LAYER Via34 ;
    RECT 63.595 0.19 65.415 9.81 ;
    LAYER Via34 ;
    RECT 72.595 0.19 74.415 9.81 ;
    LAYER Via34 ;
    RECT 81.595 0.19 83.415 9.81 ;
    LAYER Via34 ;
    RECT 90.595 0.19 92.415 9.81 ;
    LAYER Via34 ;
    RECT 100.25 0.19 107.79 9.81 ;
    LAYER Via34 ;
    RECT 124.23 0.19 127.09 9.81 ;
    LAYER Via34 ;
    RECT 129.875 0.19 130.655 9.81 ;
    LAYER Via34 ;
    RECT 132.795 0.19 133.575 9.81 ;
    LAYER Via34 ;
    RECT 135.715 0.19 136.495 9.81 ;
    LAYER Via34 ;
    RECT 138.635 0.19 139.415 9.81 ;
    LAYER Via34 ;
    RECT 147.895 0.19 148.675 9.81 ;
    LAYER Via34 ;
    RECT 150.815 0.19 151.595 9.81 ;
    LAYER Via34 ;
    RECT 153.735 0.19 154.515 9.81 ;
    LAYER Via34 ;
    RECT 156.655 0.19 157.435 9.81 ;
    LAYER Via34 ;
    RECT 159.575 0.19 160.355 9.81 ;
    LAYER Via34 ;
    RECT 162.495 0.19 163.275 9.81 ;
    LAYER Via34 ;
    RECT 165.415 0.19 166.195 9.81 ;
    LAYER Via34 ;
    RECT 174.675 0.19 175.455 9.81 ;
    LAYER Via34 ;
    RECT 177.595 0.19 178.375 9.81 ;
    LAYER Via34 ;
    RECT 180.515 0.19 181.295 9.81 ;
    LAYER Via34 ;
    RECT 183.435 0.19 184.215 9.81 ;
    LAYER Via34 ;
    RECT 186.355 0.19 187.135 9.81 ;
    LAYER Via34 ;
    RECT 189.275 0.19 190.055 9.81 ;
    LAYER Via34 ;
    RECT 192.195 0.19 192.975 9.81 ;
    LAYER Via34 ;
    RECT 201.455 0.19 202.235 9.81 ;
    LAYER Via34 ;
    RECT 204.375 0.19 205.155 9.81 ;
    LAYER Via34 ;
    RECT 207.295 0.19 208.075 9.81 ;
    LAYER Via34 ;
    RECT 210.215 0.19 210.995 9.81 ;
    LAYER Via34 ;
    RECT 213.135 0.19 213.915 9.81 ;
    LAYER Via34 ;
    RECT 216.055 0.19 216.835 9.81 ;
    LAYER Via34 ;
    RECT 218.975 0.19 219.755 9.81 ;
    LAYER Via34 ;
    RECT 228.235 0.19 229.015 9.81 ;
    LAYER Via34 ;
    RECT 231.155 0.19 231.935 9.81 ;
    LAYER Via34 ;
    RECT 234.075 0.19 234.855 9.81 ;
    LAYER Via34 ;
    RECT 236.995 0.19 237.775 9.81 ;
    LAYER Via34 ;
    RECT 239.915 0.19 240.695 9.81 ;
    LAYER Via34 ;
    RECT 242.835 0.19 243.615 9.81 ;
    LAYER Via34 ;
    RECT 245.755 0.19 246.535 9.81 ;
    LAYER Via34 ;
    RECT 255.015 0.19 255.795 9.81 ;
    LAYER Via34 ;
    RECT 257.935 0.19 258.715 9.81 ;
    LAYER Via34 ;
    RECT 260.855 0.19 261.635 9.81 ;
    LAYER Via34 ;
    RECT 263.775 0.19 264.555 9.81 ;
    LAYER Via34 ;
    RECT 266.695 0.19 267.475 9.81 ;
    LAYER Via34 ;
    RECT 269.615 0.19 270.395 9.81 ;
    LAYER Via34 ;
    RECT 272.535 0.19 273.315 9.81 ;
    LAYER Via34 ;
    RECT 281.795 0.19 282.575 9.81 ;
    LAYER Via34 ;
    RECT 284.715 0.19 285.495 9.81 ;
    LAYER Via34 ;
    RECT 287.635 0.19 288.415 9.81 ;
    LAYER Via34 ;
    RECT 290.555 0.19 291.335 9.81 ;
    LAYER Via34 ;
    RECT 293.475 0.19 294.255 9.81 ;
    LAYER Via34 ;
    RECT 296.395 0.19 297.175 9.81 ;
    LAYER Via34 ;
    RECT 299.315 0.19 300.095 9.81 ;
    LAYER Via34 ;
    RECT 308.575 0.19 309.355 9.81 ;
    LAYER Via34 ;
    RECT 311.495 0.19 312.275 9.81 ;
    LAYER Via34 ;
    RECT 314.415 0.19 315.195 9.81 ;
    LAYER Via34 ;
    RECT 317.335 0.19 318.115 9.81 ;
    LAYER Via34 ;
    RECT 320.255 0.19 321.035 9.81 ;
    LAYER Via34 ;
    RECT 323.175 0.19 323.955 9.81 ;
    LAYER Via34 ;
    RECT 326.095 0.19 326.875 9.81 ;
    LAYER Via34 ;
    RECT 335.355 0.19 336.135 9.81 ;
    LAYER Via34 ;
    RECT 338.275 0.19 339.055 9.81 ;
    LAYER Via34 ;
    RECT 341.195 0.19 341.975 9.81 ;
    LAYER Via34 ;
    RECT 344.115 0.19 344.895 9.81 ;
    LAYER Via34 ;
    RECT 358.355 23.81 367.975 24.59 ;
    LAYER Via34 ;
    RECT 358.355 47.13 367.975 48.95 ;
    LAYER Via34 ;
    RECT 358.355 54.74 367.975 56.04 ;
    LAYER Via34 ;
    RECT 358.355 58.79 367.975 60.61 ;
    LAYER Via34 ;
    RECT 358.355 70.59 367.975 72.41 ;
    LAYER Via34 ;
    RECT 358.355 78.47 367.975 79.25 ;
    LAYER Via34 ;
    RECT 358.355 86.69 367.975 87.47 ;
    LAYER Via34 ;
    RECT 358.355 90.585 367.975 91.365 ;
    LAYER Via34 ;
    RECT 358.355 97.72 367.975 99.54 ;
    LAYER Via34 ;
    RECT 358.355 109.325 367.975 111.145 ;
    LAYER Via34 ;
    RECT 358.355 113.855 367.975 115.155 ;
    LAYER Via34 ;
    RECT 358.355 120.805 367.975 122.625 ;
    LAYER Via34 ;
    RECT 358.355 125.315 367.975 127.655 ;
    LAYER Via34 ;
    RECT 0.19 24.785 9.81 25.565 ;
    LAYER Via34 ;
    RECT 0.19 39.43 9.81 43.85 ;
    LAYER Via34 ;
    RECT 0.19 56.75 9.81 63.25 ;
    LAYER Via34 ;
    RECT 0.19 77.97 9.81 78.75 ;
    LAYER Via34 ;
    RECT 0.19 88.4 9.81 89.7 ;
    LAYER Via34 ;
    RECT 0.19 97.72 9.81 99.54 ;
    LAYER Via34 ;
    RECT 0.19 109.88 9.81 112.74 ;
    LAYER Via34 ;
    RECT 0.19 120.285 9.81 123.145 ;
    LAYER Via34 ;
    RECT 23.395 166.435 24.695 176.055 ;
    LAYER Via34 ;
    RECT 27.335 166.435 28.115 176.055 ;
    LAYER Via34 ;
    RECT 38.415 166.435 46.995 176.055 ;
    LAYER Via34 ;
    RECT 57.615 166.435 66.195 176.055 ;
    LAYER Via34 ;
    RECT 76.815 166.435 85.395 176.055 ;
    LAYER Via34 ;
    RECT 95.93 166.435 98.79 176.055 ;
    LAYER Via34 ;
    RECT 102.65 166.435 106.03 176.055 ;
    LAYER Via34 ;
    RECT 111.29 166.435 114.67 176.055 ;
    LAYER Via34 ;
    RECT 119.85 166.435 122.19 176.055 ;
    LAYER Via34 ;
    RECT 127.895 166.435 129.195 176.055 ;
    LAYER Via34 ;
    RECT 131.495 166.435 134.875 176.055 ;
    LAYER Via34 ;
    RECT 137.335 166.435 140.715 176.055 ;
    LAYER Via34 ;
    RECT 142.745 166.435 144.565 176.055 ;
    LAYER Via34 ;
    RECT 146.595 166.435 149.975 176.055 ;
    LAYER Via34 ;
    RECT 152.435 166.435 155.815 176.055 ;
    LAYER Via34 ;
    RECT 158.275 166.435 161.655 176.055 ;
    LAYER Via34 ;
    RECT 164.115 166.435 167.495 176.055 ;
    LAYER Via34 ;
    RECT 169.525 166.435 171.345 176.055 ;
    LAYER Via34 ;
    RECT 173.375 166.435 176.755 176.055 ;
    LAYER Via34 ;
    RECT 179.215 166.435 182.595 176.055 ;
    LAYER Via34 ;
    RECT 185.055 166.435 188.435 176.055 ;
    LAYER Via34 ;
    RECT 190.895 166.435 194.275 176.055 ;
    LAYER Via34 ;
    RECT 196.305 166.435 198.125 176.055 ;
    LAYER Via34 ;
    RECT 200.155 166.435 203.535 176.055 ;
    LAYER Via34 ;
    RECT 205.995 166.435 209.375 176.055 ;
    LAYER Via34 ;
    RECT 211.835 166.435 215.215 176.055 ;
    LAYER Via34 ;
    RECT 217.675 166.435 221.055 176.055 ;
    LAYER Via34 ;
    RECT 223.085 166.435 224.905 176.055 ;
    LAYER Via34 ;
    RECT 226.935 166.435 230.315 176.055 ;
    LAYER Via34 ;
    RECT 232.775 166.435 236.155 176.055 ;
    LAYER Via34 ;
    RECT 238.615 166.435 241.995 176.055 ;
    LAYER Via34 ;
    RECT 244.455 166.435 247.835 176.055 ;
    LAYER Via34 ;
    RECT 249.865 166.435 251.685 176.055 ;
    LAYER Via34 ;
    RECT 253.715 166.435 257.095 176.055 ;
    LAYER Via34 ;
    RECT 259.555 166.435 262.935 176.055 ;
    LAYER Via34 ;
    RECT 265.395 166.435 268.775 176.055 ;
    LAYER Via34 ;
    RECT 271.235 166.435 274.615 176.055 ;
    LAYER Via34 ;
    RECT 276.645 166.435 278.465 176.055 ;
    LAYER Via34 ;
    RECT 280.495 166.435 283.875 176.055 ;
    LAYER Via34 ;
    RECT 286.335 166.435 289.715 176.055 ;
    LAYER Via34 ;
    RECT 292.175 166.435 295.555 176.055 ;
    LAYER Via34 ;
    RECT 298.015 166.435 301.395 176.055 ;
    LAYER Via34 ;
    RECT 303.425 166.435 305.245 176.055 ;
    LAYER Via34 ;
    RECT 307.275 166.435 310.655 176.055 ;
    LAYER Via34 ;
    RECT 313.115 166.435 316.495 176.055 ;
    LAYER Via34 ;
    RECT 318.955 166.435 322.335 176.055 ;
    LAYER Via34 ;
    RECT 324.795 166.435 328.175 176.055 ;
    LAYER Via34 ;
    RECT 330.205 166.435 332.025 176.055 ;
    LAYER Via34 ;
    RECT 334.055 166.435 337.435 176.055 ;
    LAYER Via34 ;
    RECT 339.895 166.435 343.275 176.055 ;
    LAYER Via34 ;
    RECT 344.645 166.435 344.905 176.055 ;
    LAYER Via34 ;
    RECT 23.4 10.79 24.7 20.41 ;
    LAYER Via34 ;
    RECT 31.315 10.79 34.695 20.41 ;
    LAYER Via34 ;
    RECT 41.095 10.79 42.915 20.41 ;
    LAYER Via34 ;
    RECT 50.095 10.79 51.915 20.41 ;
    LAYER Via34 ;
    RECT 59.095 10.79 60.915 20.41 ;
    LAYER Via34 ;
    RECT 68.095 10.79 69.915 20.41 ;
    LAYER Via34 ;
    RECT 77.095 10.79 78.915 20.41 ;
    LAYER Via34 ;
    RECT 86.095 10.79 87.915 20.41 ;
    LAYER Via34 ;
    RECT 95.93 10.79 98.79 20.41 ;
    LAYER Via34 ;
    RECT 114.05 10.79 121.59 20.41 ;
    LAYER Via34 ;
    RECT 127.895 10.79 129.195 20.41 ;
    LAYER Via34 ;
    RECT 131.335 10.79 132.115 20.41 ;
    LAYER Via34 ;
    RECT 134.255 10.79 135.035 20.41 ;
    LAYER Via34 ;
    RECT 137.175 10.79 137.955 20.41 ;
    LAYER Via34 ;
    RECT 140.095 10.79 140.875 20.41 ;
    LAYER Via34 ;
    RECT 143.265 10.79 144.045 20.41 ;
    LAYER Via34 ;
    RECT 146.435 10.79 147.215 20.41 ;
    LAYER Via34 ;
    RECT 149.355 10.79 150.135 20.41 ;
    LAYER Via34 ;
    RECT 152.275 10.79 153.055 20.41 ;
    LAYER Via34 ;
    RECT 155.195 10.79 155.975 20.41 ;
    LAYER Via34 ;
    RECT 158.115 10.79 158.895 20.41 ;
    LAYER Via34 ;
    RECT 161.035 10.79 161.815 20.41 ;
    LAYER Via34 ;
    RECT 163.955 10.79 164.735 20.41 ;
    LAYER Via34 ;
    RECT 166.875 10.79 167.655 20.41 ;
    LAYER Via34 ;
    RECT 170.045 10.79 170.825 20.41 ;
    LAYER Via34 ;
    RECT 173.215 10.79 173.995 20.41 ;
    LAYER Via34 ;
    RECT 176.135 10.79 176.915 20.41 ;
    LAYER Via34 ;
    RECT 179.055 10.79 179.835 20.41 ;
    LAYER Via34 ;
    RECT 181.975 10.79 182.755 20.41 ;
    LAYER Via34 ;
    RECT 184.895 10.79 185.675 20.41 ;
    LAYER Via34 ;
    RECT 187.815 10.79 188.595 20.41 ;
    LAYER Via34 ;
    RECT 190.735 10.79 191.515 20.41 ;
    LAYER Via34 ;
    RECT 193.655 10.79 194.435 20.41 ;
    LAYER Via34 ;
    RECT 196.825 10.79 197.605 20.41 ;
    LAYER Via34 ;
    RECT 199.995 10.79 200.775 20.41 ;
    LAYER Via34 ;
    RECT 202.915 10.79 203.695 20.41 ;
    LAYER Via34 ;
    RECT 205.835 10.79 206.615 20.41 ;
    LAYER Via34 ;
    RECT 208.755 10.79 209.535 20.41 ;
    LAYER Via34 ;
    RECT 211.675 10.79 212.455 20.41 ;
    LAYER Via34 ;
    RECT 214.595 10.79 215.375 20.41 ;
    LAYER Via34 ;
    RECT 217.515 10.79 218.295 20.41 ;
    LAYER Via34 ;
    RECT 220.435 10.79 221.215 20.41 ;
    LAYER Via34 ;
    RECT 223.605 10.79 224.385 20.41 ;
    LAYER Via34 ;
    RECT 226.775 10.79 227.555 20.41 ;
    LAYER Via34 ;
    RECT 229.695 10.79 230.475 20.41 ;
    LAYER Via34 ;
    RECT 232.615 10.79 233.395 20.41 ;
    LAYER Via34 ;
    RECT 235.535 10.79 236.315 20.41 ;
    LAYER Via34 ;
    RECT 238.455 10.79 239.235 20.41 ;
    LAYER Via34 ;
    RECT 241.375 10.79 242.155 20.41 ;
    LAYER Via34 ;
    RECT 244.295 10.79 245.075 20.41 ;
    LAYER Via34 ;
    RECT 247.215 10.79 247.995 20.41 ;
    LAYER Via34 ;
    RECT 250.385 10.79 251.165 20.41 ;
    LAYER Via34 ;
    RECT 253.555 10.79 254.335 20.41 ;
    LAYER Via34 ;
    RECT 256.475 10.79 257.255 20.41 ;
    LAYER Via34 ;
    RECT 259.395 10.79 260.175 20.41 ;
    LAYER Via34 ;
    RECT 262.315 10.79 263.095 20.41 ;
    LAYER Via34 ;
    RECT 265.235 10.79 266.015 20.41 ;
    LAYER Via34 ;
    RECT 268.155 10.79 268.935 20.41 ;
    LAYER Via34 ;
    RECT 271.075 10.79 271.855 20.41 ;
    LAYER Via34 ;
    RECT 273.995 10.79 274.775 20.41 ;
    LAYER Via34 ;
    RECT 277.165 10.79 277.945 20.41 ;
    LAYER Via34 ;
    RECT 280.335 10.79 281.115 20.41 ;
    LAYER Via34 ;
    RECT 283.255 10.79 284.035 20.41 ;
    LAYER Via34 ;
    RECT 286.175 10.79 286.955 20.41 ;
    LAYER Via34 ;
    RECT 289.095 10.79 289.875 20.41 ;
    LAYER Via34 ;
    RECT 292.015 10.79 292.795 20.41 ;
    LAYER Via34 ;
    RECT 294.935 10.79 295.715 20.41 ;
    LAYER Via34 ;
    RECT 297.855 10.79 298.635 20.41 ;
    LAYER Via34 ;
    RECT 300.775 10.79 301.555 20.41 ;
    LAYER Via34 ;
    RECT 303.945 10.79 304.725 20.41 ;
    LAYER Via34 ;
    RECT 307.115 10.79 307.895 20.41 ;
    LAYER Via34 ;
    RECT 310.035 10.79 310.815 20.41 ;
    LAYER Via34 ;
    RECT 312.955 10.79 313.735 20.41 ;
    LAYER Via34 ;
    RECT 315.875 10.79 316.655 20.41 ;
    LAYER Via34 ;
    RECT 318.795 10.79 319.575 20.41 ;
    LAYER Via34 ;
    RECT 321.715 10.79 322.495 20.41 ;
    LAYER Via34 ;
    RECT 324.635 10.79 325.415 20.41 ;
    LAYER Via34 ;
    RECT 327.555 10.79 328.335 20.41 ;
    LAYER Via34 ;
    RECT 330.725 10.79 331.505 20.41 ;
    LAYER Via34 ;
    RECT 333.895 10.79 334.675 20.41 ;
    LAYER Via34 ;
    RECT 336.815 10.79 337.595 20.41 ;
    LAYER Via34 ;
    RECT 339.735 10.79 340.515 20.41 ;
    LAYER Via34 ;
    RECT 342.655 10.79 343.435 20.41 ;
    LAYER Via34 ;
    RECT 347.755 25.695 357.375 26.475 ;
    LAYER Via34 ;
    RECT 347.755 42.83 357.375 44.65 ;
    LAYER Via34 ;
    RECT 347.755 49.65 357.375 51.47 ;
    LAYER Via34 ;
    RECT 347.755 68.175 357.375 69.475 ;
    LAYER Via34 ;
    RECT 347.755 73.05 357.375 73.83 ;
    LAYER Via34 ;
    RECT 347.755 79.89 357.375 80.67 ;
    LAYER Via34 ;
    RECT 347.755 88.35 357.375 89.65 ;
    LAYER Via34 ;
    RECT 347.755 96.3 357.375 97.08 ;
    LAYER Via34 ;
    RECT 347.755 100.22 357.375 101.52 ;
    LAYER Via34 ;
    RECT 347.755 117.065 357.375 119.925 ;
    LAYER Via34 ;
    RECT 347.755 134.395 357.375 136.735 ;
    LAYER Via34 ;
    RECT 347.755 137.655 357.375 139.995 ;
    LAYER Via34 ;
    RECT 347.755 140.915 357.375 143.255 ;
    LAYER Via34 ;
    RECT 347.755 144.175 357.375 146.515 ;
    LAYER Via34 ;
    RECT 347.755 147.435 357.375 149.775 ;
    LAYER Via34 ;
    RECT 347.755 150.695 357.375 153.035 ;
    LAYER Via34 ;
    RECT 347.755 153.955 357.375 156.295 ;
    LAYER Via34 ;
    RECT 347.755 157.215 357.375 159.555 ;
    LAYER Via34 ;
    RECT 347.755 161.285 357.375 163.625 ;
    LAYER Via34 ;
    RECT 10.79 30.88 20.41 35.3 ;
    LAYER Via34 ;
    RECT 10.79 46.41 20.41 49.27 ;
    LAYER Via34 ;
    RECT 10.79 64.2 20.41 67.58 ;
    LAYER Via34 ;
    RECT 10.79 72.995 20.41 73.775 ;
    LAYER Via34 ;
    RECT 10.79 79.89 20.41 80.67 ;
    LAYER Via34 ;
    RECT 10.79 86.7 20.41 87.48 ;
    LAYER Via34 ;
    RECT 10.79 96.015 20.41 96.795 ;
    LAYER Via34 ;
    RECT 10.79 105.09 20.41 107.95 ;
    LAYER Via34 ;
    RECT 10.79 124.725 20.41 127.585 ;
    END
  #BEGINEXT "VSI SIGNATURE 1.0"
    #CREATOR "Artisan Components, Inc." ;
    #DATE "2001-05-17" ;
    #REVISION "1.0" ;
    #ENDEXT
  END rom_512x16A

MACRO pllclk
  CLASS BLOCK ;
  FOREIGN pllclk 0 0 ;
  ORIGIN 0 0 ;
  SIZE 300.00 BY 280.00 ;
  SYMMETRY X Y R90 ;
  PIN ibias
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT   0.00 185.00   0.30 186.00 ;
      END
    END ibias
  PIN refclk
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT   0.00 145.00   0.30 146.00 ;
      END
    END refclk
  PIN vcop
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.528 ;
    ANTENNAPARTIALMETALAREA 0.5819 LAYER Metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT   0.00 105.00   0.30 106.00 ;
      END
    END vcop
  PIN vcom
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.528 ;
    ANTENNAPARTIALMETALAREA 0.5819 LAYER Metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT   0.00  65.00   0.30  66.00 ;
      END
    END vcom
  PIN reset
    DIRECTION INPUT ;
    AntennaGateArea  0.792 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT   0.00  25.00   0.30  26.00 ;
      END
    END reset
  PIN clk1x
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.528 ;
    ANTENNAPARTIALMETALAREA 0.5819 LAYER Metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 299.30 185.00 300.00 186.00 ;
      END
    END clk1x
  PIN clk2x
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.528 ;
    ANTENNAPARTIALMETALAREA 0.5819 LAYER Metal1 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8143 LAYER Metal1 ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
      RECT 299.30 145.00 300.00 146.00 ;
      END
    END clk2x
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
#     SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.00 235.00 2.00 245.00 ;
      LAYER Metal3 ;
      RECT 0.00 235.00 2.00 245.00 ;
      END
    END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
#     SHAPE RING ;
    PORT
      LAYER Metal5 ;
      RECT 0.00   5.00 2.00  15.00 ;
      LAYER Metal3 ;
      RECT 0.00   5.00 2.00  15.00 ;
      END
    END gnd!
  OBS
    LAYER OVERLAP ;
    RECT 0.00 0.00 300.00 280.00 ;
    LAYER Metal1 ;
    RECT 0.30 0.00 299.30 280.00 ;
    LAYER Metal2 ;
    RECT 0.30 0.00 299.30 280.00 ;
    LAYER Metal3 ;
    RECT 0.30 0.00 299.30 280.00 ;
    LAYER Metal4 ;
    RECT 0.30 0.00 299.30 280.00 ;
    LAYER Metal5 ;
    RECT 0.30 0.00 299.30 280.00 ;
    LAYER Metal6 ;
    RECT 0.30 0.00 299.30 280.00 ;
    END
  #BEGINEXT "Created By:"
    #CREATOR "Cadence Design Systems, Inc." ;
    #DATE "2001-04-27" ;
    #REVISION "1.0" ;
    #ENDEXT
  END pllclk

MACRO ANTENNA
  CLASS CORE ANTENNACELL ;
  FOREIGN INVX1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.32 BY 5.04 ;
  SYMMETRY X Y ;
  SITE tsm3site ;

  PIN A
  DIRECTION INPUT ;
  ANTENNADIFFAREA 0.7845 ;
     PORT
      LAYER Metal1 ;
      RECT 1.065 2.37 1.18 3.56 ;
      RECT 0.835 1.35 1.065 3.56 ;
      RECT 0.8 2.37 0.835 3.56 ;
     END
  END A

  PIN VSS
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 -0.4 1.32 0.4 ;
      RECT 0.18 -0.4 0.52 0.575 ;
      RECT 0 -0.4 0.18 0.4 ;
     END
  END VSS

  PIN VDD
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
     PORT
      LAYER Metal1 ;
      RECT 0.52 4.64 1.32 5.44 ;
      RECT 0.18 4.465 0.52 5.44 ;
      RECT 0 4.64 0.18 5.44 ;
     END
  END VDD
END ANTENNA

END LIBRARY
